PK
     T\:�b��N  �N     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8"],"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9"],"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5"],"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2"],"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3"],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7"],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9"],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13"],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12"],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_4":[],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_5":[],"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_6":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_0":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_1":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_4":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_6":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_10":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_11":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2"],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_14":[],"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_15":[]},"pin_to_color":{"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0":"#010067","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1":"#9E008E","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2":"#0E4CA1","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3":"#FFE502","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4":"#005F39","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0":"#95003A","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1":"#9E008E","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2":"#FF937E","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3":"#001544","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_4":"#000000","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_5":"#000000","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_6":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_0":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_1":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2":"#FFE502","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3":"#005F39","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_4":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5":"#0E4CA1","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_6":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7":"#95003A","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8":"#010067","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9":"#9E008E","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_10":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_11":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12":"#001544","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13":"#FF937E","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_14":"#000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_15":"#000000"},"pin_to_state":{"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0":"neutral","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1":"neutral","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2":"neutral","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3":"neutral","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_4":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_5":"neutral","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_6":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_0":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_1":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_4":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_6":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_10":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_11":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_14":"neutral","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_15":"neutral"},"next_color_idx":8,"wires_placed_in_order":[["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8"],["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9"],["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5"],["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3"],["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4"],["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7"],["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1"],["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13"],["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8"]]],[[],[["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9"]]],[[],[["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5"]]],[[],[["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3"]]],[[],[["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4"]]],[[],[["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7"]]],[[],[["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1"]]],[[],[["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13"]]],[[],[["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0":"0000000000000000","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1":"0000000000000001","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2":"0000000000000002","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3":"0000000000000003","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4":"0000000000000004","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0":"0000000000000005","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1":"0000000000000001","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2":"0000000000000006","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3":"0000000000000007","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_4":"_","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_5":"_","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_6":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_0":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_1":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2":"0000000000000003","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3":"0000000000000004","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_4":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5":"0000000000000002","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_6":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7":"0000000000000005","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8":"0000000000000000","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9":"0000000000000001","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_10":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_11":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12":"0000000000000007","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13":"0000000000000006","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_14":"_","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_15":"_"},"component_id_to_pins":{"03ba13d2-1393-4316-9b38-bc1aad520043":["0","1","2","3","4"],"4144bdea-100b-4a9a-af20-60ffe64f4a21":["0","1","2","3","4","5","6"],"efee3ff0-6a5f-4fee-8269-fdead77a32d9":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8"],"0000000000000001":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9","pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1"],"0000000000000002":["pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5"],"0000000000000003":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3"],"0000000000000004":["pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3","pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4"],"0000000000000005":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7"],"0000000000000006":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13"],"0000000000000007":["pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3","pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000006":"Net 6","0000000000000007":"Net 7"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[1050.2784955,166.18519100000003],"typeId":"63e1dcb4-70d2-41a3-ab14-cb1f0167e7ff","componentVersion":1,"instanceId":"03ba13d2-1393-4316-9b38-bc1aad520043","orientation":"up","circleData":[[587.5,125],[586.6165,142.664],[585.733,162.9770000000001],[588.3834999999999,183.29150000000004],[587.5,201.83900000000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1081.7697309999999,418.41351499999996],"typeId":"04ca8eb3-fe95-4482-8406-ce523551a7a7","componentVersion":1,"instanceId":"4144bdea-100b-4a9a-af20-60ffe64f4a21","orientation":"up","circleData":[[1022.5,319.99999999999994],[1022.1952884999998,335.1809015],[1022.4904839999999,350.85205099999996],[1022.150623,366.48518149999995],[1022.4904839999999,381.778448],[1021.8107605,397.41152],[1022.4904839999999,413.04464899999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[774.6732715,453.086372],"typeId":"999f3859-f3cf-40a6-9c15-be46b91481ac","componentVersion":1,"instanceId":"efee3ff0-6a5f-4fee-8269-fdead77a32d9","orientation":"up","circleData":[[707.5,395],[707.5,410],[707.5,425],[707.5,440],[707.5,455],[707.5,470],[707.5,485],[707.5,500],[842.5,500],[842.5,485],[842.5,470],[842.5,455],[842.5,440],[842.5,425],[842.5,410],[842.5,395]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"42.07524","left":"568.13137","width":"964.29425","height":"521.99541","x":"568.13137","y":"42.07524"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8\",\"rawStartPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_0\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_125.0000000000\\\",\\\"542.5000000000_125.0000000000\\\",\\\"542.5000000000_335.0000000000\\\",\\\"887.5000000000_335.0000000000\\\",\\\"887.5000000000_500.0000000000\\\",\\\"842.5000000000_500.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9\",\"rawStartPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_1\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"586.6165000000_142.6640000000\\\",\\\"572.0582500000_142.6640000000\\\",\\\"572.0582500000_140.0000000000\\\",\\\"527.5000000000_140.0000000000\\\",\\\"527.5000000000_305.0000000000\\\",\\\"902.5000000000_305.0000000000\\\",\\\"902.5000000000_485.0000000000\\\",\\\"842.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9\",\"rawStartPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_1\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.1952885000_335.1809015000\\\",\\\"1007.3476442500_335.1809015000\\\",\\\"1007.3476442500_335.0000000000\\\",\\\"902.5000000000_335.0000000000\\\",\\\"902.5000000000_485.0000000000\\\",\\\"842.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5\",\"rawStartPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_2\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"585.7330000000_162.9770000000\\\",\\\"571.6165000000_162.9770000000\\\",\\\"571.6165000000_170.0000000000\\\",\\\"512.5000000000_170.0000000000\\\",\\\"512.5000000000_470.0000000000\\\",\\\"707.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2\",\"rawStartPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_3\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"588.3835000000_183.2915000000\\\",\\\"572.9417500000_183.2915000000\\\",\\\"572.9417500000_185.0000000000\\\",\\\"497.5000000000_185.0000000000\\\",\\\"497.5000000000_425.0000000000\\\",\\\"707.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3\",\"rawStartPinId\":\"pin-type-component_03ba13d2-1393-4316-9b38-bc1aad520043_4\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_201.8390000000\\\",\\\"557.5000000000_201.8390000000\\\",\\\"557.5000000000_440.0000000000\\\",\\\"707.5000000000_440.0000000000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7\",\"rawStartPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_0\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_320.0000000000\\\",\\\"992.5000000000_320.0000000000\\\",\\\"992.5000000000_297.5000000000\\\",\\\"1180.0000000000_297.5000000000\\\",\\\"1180.0000000000_575.0000000000\\\",\\\"670.0000000000_575.0000000000\\\",\\\"670.0000000000_500.0000000000\\\",\\\"707.5000000000_500.0000000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13\",\"rawStartPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_2\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.4904840000_350.8520510000\\\",\\\"1007.4952420000_350.8520510000\\\",\\\"1007.4952420000_350.0000000000\\\",\\\"872.5000000000_350.0000000000\\\",\\\"872.5000000000_425.0000000000\\\",\\\"842.5000000000_425.0000000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3\",\"endPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12\",\"rawStartPinId\":\"pin-type-component_4144bdea-100b-4a9a-af20-60ffe64f4a21_3\",\"rawEndPinId\":\"pin-type-component_efee3ff0-6a5f-4fee-8269-fdead77a32d9_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.1506230000_366.4851815000\\\",\\\"992.5000000000_366.4851815000\\\",\\\"992.5000000000_440.0000000000\\\",\\\"842.5000000000_440.0000000000\\\"]}\"}"],"projectDescription":""}PK
     T\               jsons/PK
     T\�#��(  (     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"MAX7219 8x32 LED Matrix","category":["User Defined"],"id":"63e1dcb4-70d2-41a3-ab14-cb1f0167e7ff","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"41d41cfa-55db-4eb2-805f-824b346b9186.png","iconPic":"2dd0ce04-414d-4887-acda-26c206c9abda.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"62.95295","numDisplayRows":"15.21466","pins":[{"uniquePinIdString":"0","positionMil":"62.45753,1035.30094","isAnchorPin":true,"label":"Vcc"},{"uniquePinIdString":"1","positionMil":"56.56753,917.54094","isAnchorPin":false,"label":"Gnd"},{"uniquePinIdString":"2","positionMil":"50.67753,782.12094","isAnchorPin":false,"label":"Din"},{"uniquePinIdString":"3","positionMil":"68.34753,646.69094","isAnchorPin":false,"label":"CS"},{"uniquePinIdString":"4","positionMil":"62.45753,523.04094","isAnchorPin":false,"label":"CLK"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"SCD30","category":["User Defined"],"id":"04ca8eb3-fe95-4482-8406-ce523551a7a7","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d10c801-e2f1-4174-9a9c-587482dea60d.png","iconPic":"05c4396c-27e7-4cac-a4cc-0e5db7270844.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"9.05512","numDisplayRows":"14.17323","pins":[{"uniquePinIdString":"0","positionMil":"57.62446,1364.75160","isAnchorPin":true,"label":"Vin"},{"uniquePinIdString":"1","positionMil":"55.59305,1263.54559","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"57.56102,1159.07126","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"3","positionMil":"55.29528,1054.85039","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"4","positionMil":"57.56102,952.89528","isAnchorPin":false,"label":"RDY"},{"uniquePinIdString":"5","positionMil":"53.02953,848.67480","isAnchorPin":false,"label":"PWM"},{"uniquePinIdString":"6","positionMil":"57.56102,744.45394","isAnchorPin":false,"label":"SEL"}],"pinType":"wired"},"properties":[],"hasComponentImageSvg":false,"componentImageSvgUrl":""},{"subtypeName":"Wemos D1 Mini","category":["User Defined"],"id":"999f3859-f3cf-40a6-9c15-be46b91481ac","userDefined":true,"subtypeDescription":"","subtypePic":"f814d8c7-8d80-4469-af20-bcf736e1bcac.png","pinInfo":{"numDisplayCols":"10.07874","numDisplayRows":"13.46457","pins":[{"uniquePinIdString":"0","positionMil":"56.11519,1060.47098","isAnchorPin":true,"label":"RST"},{"uniquePinIdString":"1","positionMil":"56.11519,960.47098","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"2","positionMil":"56.11519,860.47098","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"3","positionMil":"56.11519,760.47098","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"4","positionMil":"56.11519,660.47098","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"5","positionMil":"56.11519,560.47098","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"6","positionMil":"56.11519,460.47098","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"7","positionMil":"56.11519,360.47098","isAnchorPin":false,"label":"3V3"},{"uniquePinIdString":"8","positionMil":"956.11519,360.47098","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"9","positionMil":"956.11519,460.47098","isAnchorPin":false,"label":"G"},{"uniquePinIdString":"10","positionMil":"956.11519,560.47098","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"11","positionMil":"956.11519,660.47098","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"12","positionMil":"956.11519,760.47098","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"13","positionMil":"956.11519,860.47098","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"14","positionMil":"956.11519,960.47098","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"15","positionMil":"956.11519,1060.47098","isAnchorPin":false,"label":"TX"}],"pinType":"wired"},"properties":[],"iconPic":"858a2a89-b1fb-4d30-9067-568b89f7eae7.png","componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     T\               images/PK
     T\ѥ� �� �� /   images/41d41cfa-55db-4eb2-805f-824b346b9186.png�PNG

   IHDR  �   �   +�   	pHYs  �  ��+  ��IDATx���w�,E��_={�^1��A$�d$	�E�����EQ�(b�0���$
�I�9KF0�{=gO�>O�O��5�ӽ�����y��Z�»V�Z5Y�u�?4~��{�p�	3�g0�M�'&&�<�'}۪�ү���fϞ���<������ÚN������x0Ř����-��瓓����|���{�h.�QM;α}�V']��?6z�_�_5M�OK��'���_#WD��K��ճf��_��k���>�=S?��ćs�&~Q
|h�����q�QW��8T�H�%����x22��U#�-�b��S��<>�ᩥ���:�t���O lduu�C������9Vͼy튡�^:�~�o������?;��g��Bgj<���bZ.j��-GUn��H��m쐊ŝa+��</vM3^��O��Rн�Ђ�gb&
"h=���CJjRf�� i�����������8��,Aԁh�aӊ��GE$ݮ�~��>�Cz��`�q��W㜡�V{�s���h->���`��z��AEd���	��6s��� �����9֔�_��X�M�ʳ����������+�<hZA�9y\��E�iT�n��v�d�77O�H£/@s?�d���M��4g��{���*]�{$�(��]Դ�s��������O� ���C1=S�al�zT��Կ���s�Fb|��5 ��[*̾z�5�JOW���I'�J��sW'҉����v��,a>��m�?��bv)S���?C����*�/�P���]�^M���HC��b���4�wgGB��2I���^\�W=�"�:��'�/�%��T�=�G=����kN�ł#0��DK�����4�B{��b����'�=��x��ȦT������ot�%�|�?�����=O0����'����h�_C�be�^a>�V,�g5ڑK��cl�r����ixQ�����X_~�8~]ъ��$�S�m�")�U�d$�z�!AT&��z�0��Hw�[�c�C)k���E��FP���-p�>����5j�ii�C�ҡ����f_N�d�)�Z���{�q�q�fs������/��9���οZS=Y :{Aj4s3�cy��[WDmك���_�/�Ն�6{q!�H�b��BH�QDt.���<܅�SP%Q�����p��ߢۖ�$�O<�0�;�~h{/S�򍍜�;-��WK���}�5o
�N�9�lg�̀�^����Y@�����FU^����ֆ��@8>cD"��l�ӳp]<�h'R��"��,��F
x�)k�">GݶY ��Lkod%J�����G�,�lY�y����3�^������Х����Z�#�����:#�6�I�J�^���{��K (���D[�����5��2���a��R���Pä��pD���o6#��� �y&���iS�y'v��|vޗ��}`ۻ�(���Ty�8��E�2e�A���~{'RhK/�W3��\���#��</��>�^�*�Kb�H��V
1+[��PZT�=��A����ÈV�3B:��<i%�����̇Z#�n_��(CU�A?�m���Hx-kd�����Wa����Gh� ���m���.���12��2����ğ���P�;�����qZ,�{�`�|f�G�P��o��)c�"�f��
�GT$��m�XB^KND�</��c�������{��Z6Kx��T��fw���طG�Ռ������� "C̩I�ؒ���#����V���an�3��&���՞�?h�QbV�>�e��6GVy���Vܮ(N4N6�sD�h�_U9�g��79]S�s�u�D["��խ�ld�Й���S�WF��P��{��yd�[��"�3��ѸT����Ԉ�%�03���衿�wv�9"�."� ��i\E"h͌�7GM*�Z�3WG.�?i+h��#���ż�am�8�VX�ht�W��������r]��9c����(eR�J��?�̙v�l,����,�vQ����gh�a�|�x�;���@�~�},ڃѝ϶�1��[
$2̵�^��J���u`�����;i21�=j#�L�?���8fW7!Ř�իiO��Eĕ������u5�#5�/�4�PTRT;�\J�l����5��^RG�������u�+f3b�$N�/5W؂�3���{���|��f뙀E�I?)���gɃ�>�}�FA�Ա���:����q�"��je��Q��aG!u���V�x��3r,!����3C��ͯ��Ѐed�"O���gw���Y�;�c��s�PT��i��xL�(\��1��[�8~�֦:��c�qA��)���qe����F�K�6�U6�Sѝ�2MM��.V�,W�:�6������y�.V�C�d�X�	o_ё�����c��x�s��l #T�po��*�Ҩa{��H�Q�9�j4R5ș?O��O�f���˄m�?���A�%ư_�m�t^ө�5��H�c�S9R�6HM��B4G��iƸ_�J�TywBz�
9u=r:�����/e17��H�LyS�k��S|���>�I�G�9�����ڊ�n��0�f<0�)�`�dM����D;?���Կ�q������S�����Qh�O�I�>Ex�_�ۀ6��z��C��B5`��Fa��Z�M����q�e0�t���{`bc������`����c@Y��iuiR�m���+�)H��k�1z��:�=5����0o@I�����#���iL�{��X`��矟��O���׿>��S�.��=\�I2=>+X�5��/�0���������/�K���c'�4�-ea����E��7����_�9�~�駭%�����VK�>���/]p����z�XUW�ǰ�D6�5����/\h��^���?���>�����ߢ�̑�t���j3<�'�x��S���@��ς���_�b��F?���?XJ<�c:�T�|��a�9���t+*�<�{P��k�)�K��_V�%�]�	��g�yFA�❡wd�����*��ЇY����qfB�4�(y�(CҳHC2rq�z�u_T��gX�ӳ�5�=3x˂�ԣm�v-PL��w�y�Q5��	�z�ˎA�*�rʍ �g�t�H�Í�<�H;
�M�(���c��>�s^Ā}�Q�t"�1��:ƷX���c0	#�g��'�����z4�u�if��->,x���R���P���:�6�{���R��v�0�WPU���.�$�������9+�$�(�1x�Lb�����9"�C�/��t��vo/��i��=-.�D0lh��ax�k���z�lχ����u4�Q�H7�c=]�iLIb��7M4�O�	|�K�d>f�#p��A=M 8�""`�0I<2�aٴܮ˛M�� ;S`eŐ����ɍ��`��
��$&
�@�EYDJ�7ҳ�d�X����$�W|`��$��؃n�)�k��$2G9�x�oT9�F�b�4�l�v��*Z{���P٧gԻ�=r�o���P0	��8Q�(��0줍��v���]��a>�~o�u�D?�-(�_��
FΗ�	B��m�R�a��n��������0�j�����ۿ�U�Z|��+#��{��⊳�>����z����	�	!�9a�[n��v�m����#3PA����N���~w�e��+r�Z�.a��$����!=��l �B���+�?��_��Wiȝ2J�G����P���C�_b�%0���O����/��l'��4�&K�P�b�-��W��կ~���n��RK������;�.�� x�?):�R�r��Yf�e5�^{m�F 鍊n:묳~���^w�u�\�~���@ƕVZ����j��[��D��y晐����gq'�fH�n~�Ou#{|��B�W��/{�� 8�E��{�ЄW`�&���~�����z1��W_�)�.�R�'X�5��o~�,$�]��yC�0�]w�u��6C��P+���׿������4�����:Q#_~���׼�50+�<�o�!�s��Nq{���@�+��?4�|�ͷ�b�e�]�Y�þ��[��_^~��t�B>^O����4\,L�m�Ѫ���t�YVx���Pp̾����l�o�++w�����������[�����N@�*�_q�_���n��6p;ɗp;�������HN� ��k�	��/��Q��D�>a��/�7	�m�BH�Az��mP;(I�A�#P5MN)�o9�h���$#�(V%I't�/z�B�k�������]0=��{Y(���뮻��:����G�ð���+7��OK1DXy�aHx�%�� 	�-g�qK���b�܍s
^��Ej0:��~YY�`HL��k=��.�����	% &Xʭ��z�M6lI^}��ػ�O?�a��1h��c�V���9z����p���^J�/��l�j��E�:���yF��v[:G`�	/�X�-���c�<�j]?V7�Y�ՊV�E(vn��	݅� �p��-C��v�)-M�X ���w�q�u�Y�ΡԾ뮻�\��Dt�@��s6
XD�=}���7Bm�5���(7���˴z���-p;rL���?d�X::�硉��f�$X
�n���\���Ub�Xp�#� V�;�,%���$�hH9�V�3M�,+�+M���w�8�0�w�Vؤi��C[�������%��Q���$�c`�@��N;��Q/�����SO��Y|R�T������?�_��*��Moz��_�Z���+7�	�g�;�8���s�@�e!�a�}�]c�5 n�ˀ|�8��o~3������R��N I-P�MB��v�m�=��?B��x�F~Џo������x���H�K?��[���v��T�C���u�{���#�8B
ќ�Q|>@H���wn��ƀ	xk�S��6�w���¶�9?��4��M�W���z�a��!�����{�t�I��[nI3n�饗~�[��@yE��(��7H��5����?G�J�th� �B�1�����p˒K.�#S�'V���~���F���~�3X1���9j�Ȉ�>�V��!�Ⲳ@^V�x�1���=�K�v�yg(�,�l��s� ����O~��]O`���;����G?
Ld����E'0˽�{�����/���7�ͯ�֖$aaYJh�r�V�&�utr*B�O��SHM����g��L%�`�kA���mo�&?��O1)۪�ğx��b��Kln�C�����YM�0�6����n�S�!���7��W8@?aFx2,"|�G�x�3dE�)�C;A,=[��I8��d�UV��A�~8@�b�O����ר�	b�u�C,3��AXq�9�����?]!��c`�%~c������!1��<�zq�x/��e�]�cp&®M$u�yӰ���N8��{�#�И;Jl��w��M4)L�Vp;l� 
�$B&�'��Z��}/��袋Xkc�v��2��z��t{��X%x�I�2��P0��'�Yn��f!��E�z��M�B50�cC�Í8���~;f��}�Qi~����^� `��	�4"��>�����"�p�l�,����~Kċ����qf���c�v #�c=J�ۧR��<�:k�X�gX\����j��=~��&���1���N��\^��D�n��6���|g�9�=�S�&#���nCj3����h6�H�A	�۫�m]�A���!��;K(%��j���	��@�.V������z�|h�qФ��/��?� ����<�B�(̝a����Sc�x ��7�x#���/�*���i4�� N36�M'1�	��%�\����b)���\����a��k_�^pJR��r�Fh���}�{_�җ�<ǹ�9�= q?�O�Q�'U(���/����Zx�cүc
(ك>�y�_뼽�������^{�}�Cw�}���zH�=�C=��C��K�	���o5͇k��_� ��?�	�vN�
>�J�%&�����	�����O��X5�� `տR%�
����x��A��\�-e���&i=Q�v�aLY��aW�2�E�a�<���л~P�V��c�9��0�CN"����n����H��Z��G`1U���E
V����_Q+G��|�Za�X�EY�a�uo̟���B`z�-,�e�:Eb��x`���=U�g�,�Q=I�c�\~�翨Z,��x(j6ML��@X0��(J�x��Y�� (A/P�)j1�	?�~T1@��y�Q(���! �2�t�AqV/�:�y/�@���[oU����Z�c��`�o~�J�d���4�u�]�	����y�0�]�Ğ�A���X�,k]+�n��_�o�ט6Ǆ�_��w��]�JVSL����Ha��������+�6I�c������/�G5��ZЀ`���sΩG��6O��&>|�n��8��Q��|�����g?��&���=���b�a;8�[>��?��1�:4�i��n<�4}�3�Qe*o�:�3���c
W�p�8J�" ibا�~�Oьm1Q���4� [����Zj����o?,5�<�a�q�.��n���>����dj�g@� X��Y�CU������G?��6W%_��VnW@�LT�N��q]��[�c�b�_�1H������`a��Ȣ���b����v�8J�5D�@I`���)7���NS�1�%W�a�5F�E+5��]�z���61zz*�
T"J��Y�o��h�ݧ-@|�;�K��~M2��r<d��X%$1����	��	�$#��Z�����h�a~%�T�h�M9R�b��!o��:�B���+����l�RƐ,7��,b:m���@�'<44ᷩ9���D�'^�P|�s���2E�nVIs�������O~�!9�K"l'�����p6�Eo�f̚Jٰy��oX���I!p��i���+8�G�!AM�CYf�4*WfqVQ:�~��e`z-��UG}�_S����(���`5���p[
���h��~��:� @/�!�����1�O}�St{�i�����;���L�<��'�*��J л0��篽�Z�kW�2�D�t4����%V@�̹�]�z�3�t,x��'��k�y����&�GiA #��U9�j��1ƨ'��,��u)Ԗ��D�N� �l϶
uvʪ�%@<�q�VXjc�?A)�� T�7�͍����BHt�Eiv���*�{I����N�]��>��hm�܎-Q�{�G�6�yC��4_�H�Caڷ�����y��Sw1�	 �x�����1SV����϶'�ơ�	����s�=����ƃc��/��t�M)s�s Rc96� ��馛������ѝɦT���l��?�&Y��0���j�C@`ej�M�Պ+e�Ɵ�%`�3�<s�)�@"�:2ș�]S�ϑq~�w��K����w_z������+Ի���<$�(H��O���=����۱p\p��%X6���3`�#ܟFw5��",(�_W���P����7�{���Q8�py��b�YY�?�sUa���@ְ��m����f S�++ǆ9>X#���2\���[���7��C�)��ꪫ~��G}������[�O2�%�\��a�rX_��$�R�W��	�ůĨ 3�)^�yUjǏ�i�q� 5���A��.�/F�!@��_Zw������{�����{��^�M���q�򕯀dR��c��I���|�Y��h�(�ʲ������;�5_$�������l��,饀c���믟�|�Wg85�������E�}���ױ�6�ғ�
,
��H��$B%RF�B|�@�0�v���V�܎� 7bO�cDK�_�P0!6����|��o����l�~�r����s�94aj������vq�'n�/�S�y�S<F���_W�\����d� ���������p�?��x�ꫯ��K
mR�`�֒i�p �e��Q� �����|���_�C�]S��aIxؙı��C�!��{H���M���1��E4�h�1���^{�z뭿�կ&� q��=<����W�� mMV��� ��^}��1�t~��ے�(g;�_�%c�x��A��X��_��W�{���?���u[�"xɟ��w��5�1m>�X:�\ 8���#��P�G���m
1�?�O�������s�u�]׵.2������
�&r�>d��~���o��n���/���p����(b�[D�1��&t΋�v��-����O�u}~�N0T���*Ri�z�0�ox���K|$��qQ�Ë�{��@�Q�u-4#���UWik�KN��a�0�����1�ڏ߰�w�}w݄����/���;���y�x ]�Px^#�,�I����*�̇���������ʅ��� �������OF�/�������_~�1\�K�wA��b�-�p���>t�-@Ư����?�L��K�f ��.!c��V�Cՠǰs�KP�����]��;��n�l�X�6���)�b4�V[mE��-�� �����h��>[n��������d��	z�[ߊ�9���q=~X�U�4Ѿe����t�=<X�޵.<�n���H�zV��ż�΋n�s8G'DS0��Oh�:N�anꆞr�w�e`�QG���L_��!�Pt���ڦ�[���?�\v�e�\�yr�^�b<�p�n*������;��3���֓N@�!J���m�4L9�_i����ң�>���qO�zl�wɼ�E/J�Y�	a�<&h���LW
e�R�&��D��9);�Jp�}K����^xa�geO=��"<Z�����+���z�=M9$�>��#x �9��"<�W/;v�8�6�l�.Rȸ ��+c�|}��uG���2���=0��	����j��N,�����D+��B�UMm"�XmU +Űwx8p;0 Q�l�CHs�k�e�!���o��bi[(F�>E�W\q��\����!���W����m�������>���;��a��p��yLg����3���omUȓ�4(A�^:��%�B,�R�c
G��i����7��o��6��.�&�l���L����h,E|h�Yt�E�Z���2l_Bp0�Yg�e�Y�x����Yg�7��;�,ꦉ\)G�5#]p�
�F���a9�qw0u,���#$-+����Z�d�rqp"����9�Ѧ��3�:@�u�n�Ȯ)��,��r^�0'2��W�0��'f;�c`GbZ%���|���.Y/�@Q�Q/\�\��;e�ȩ�!�	���O>�����o|#]���ix0���
֡ȯ'�Y��Apx�4�w�5~��O;�4^p�]u[K�'�!��=f�O2Br��6r���U�g�i<�w�	�O�Z�򱢉\�t�W��8�::�iZ=��C����/��$�|�=�P���|C h&�����i!2�p\5�w�>��'��á�T�I�Qd�,�)���,+.���J��<� �%�	�[|��$5�"}�Ρ� ��㰴O%!J�m�3��.R[����=nG�<��$e	�ӹ�o����8����)Zٵ;ʓ�#���?ߢԣ
��Y��SNQd!���h���[o�#���:Ds�&d<w�q.��3�Ǝ?5���){b]zr*ם�[�.Ŀ�⋟y��Ѡ6�x�[ނO"�߯ �(z�� J���w����i�.� ����T��+5DI���'c�&r��6}��z�Ǔ)�D����{�����9�n7�Y���p{�~�h�� �O��x�@Xe�׆���w_��?S��-����뜵�_�"6�xc��h�/*���k���cL�[C#�^�=���LQl�|�M7Ŧ�g	i\�"(�̀��c)Qj�a�A#!����F��:�J�a�y~��7_v�e1E�3js��*����M��AO��;x�?�����y �)��?*o���h7<�*nC"��ȿVR)�{�mb ��
�d��y�]vQ����;��:����y�I'�N������C��{0�t�n"��t�����F]t�E�[��a��eU��8�:\����P����>�h�N���&�S�-e�M�T:�������nV�>8��x�D�OtH���f��v�mL�����ONḂ�ӻ[�Ч��)F�^��*���*u�GUٮ8���C\�aH����*3 l�g���L�z�n|^���7,D�����d�]w��pw��6��R��t����c4��g4�2zE��-��cf�0.JG����
�8p?����a����qMŐ{8n�=z'��&��2�0ͧr��A�L5C���|�UWy���XYL�l�}©�"�po���ח�^b�a�e��m��&�w�(�֢
Ј۝����+ Qb����~h�s~��P���k��+�TfN
e�f[F'&R����P����!���bGI�s�9E\&��	�=5`1u7����#�+dn視��Yc�5���R0���e� O�f�u���w������J+��Gy�ѫ�#���^��AN�t3�=�v!)*W{����5�B���>R�=�����ۙ$�z	�]��h��=�E�\V�Y8>6}��zi���ד�v+�6��i���>@|t����-hW�p��E�+�Yg�Dy+I=�Cɰz�<;+2�zw���v��k��6�y��W_}ut��Kd��	TXKk���a�<|��K��[ƶa.�+V������e��қۋa��K�I�c5pU�4
���<���H�N�$X���m5HR�@�W��w�}��\�՝[Gc����Fv�s�aZ�}�4�n���p�ܵ���|VN.��v�7^�򗿜iz��;��9�iį���rZ���1��&��Q�MYY{�����v��>�9�>e���l��j��=𾡷e�F)P���į�ӟ��e��P�`�ȝ��7˻`Th(Fu�)��.}F�VXa�pv>{H���h�{9��93A�b����)�̐�m�Z[(��Q���2�"��YgK։�(�V�NJ���w�E��?����Bn����h�\�B�/���Y�g�y��"q�-���Ǽ�asT�}��_�S�c=��`ڕU3�Dp�n���X�$�~���^p�]�o5��UC�z�!�����h��ΓG{fa�\��:[�o��'�p¬|uq=	���F�ñxNk�t&��`��c���Yd0Mt�Ro�h��B �N�#a�!r��⋳�QètD��Q�Ԡ(�EV��}f�i�k�m���7r�Z�K��_��BFF�Ã̶��V�uG;�'�Tp�$�#�p��;���;�Z�h���c�g�����$eBCpV��[o�
|�M�c%��Ԗp�إ���]�m��a�6��������ߣ3�A�jW�ǝ�8kj�Wۋ�1hk�8f�3�!&�t�ϭ�D�-2�N�C�);�3}�b��x�� �Ql7k$���'�<��"qζUu���u�]��ɵ@��4����g܏
L��j`V;�M<#adج,>ܞF/۩B0fk�%��'�mz�l+���~Y|$��_5��� q߾���p���C�������4����ъ�Rz��."��Z�	�t�Ǫ��؆�8���і�X95��#Lx�5׌�v.G�������&g�Z]��c_��p3^d������o�E5�z)�fH�ՔJD����.�NA
�.,ӵJœj������D�;�/���6f��M���&�B����Al*%��SHE���\���w�L��1~�ID�h��O(��Z4w]z5OS�-n������i�6�O+�A��OBpG&�� �&5o~��r�M(S�rQ|�4�N���S��W[.�����?�����C �$� Z�qX��0��i �]}��iԧ��u+�|�͗�yЮ9F��WR�L��jD���@yW`�G���ȫ栈�U]�#�p�<��w��mN�h��6?��괌0� _��zc9 S}�����dd�L�R$�␉\{��Q9{J���U"cv(ە��"���e�R�dlV��e�\!�������oH04z/]�W9��/F�@�����--�8�#���H�E�H%�bn��p�53��mH�����v)I��/x�9ִ10�_4�;�Xג�E�C�T��u��
d�����ÖP�:D����%���^�^�ű`�}�u@�}|(��|�VS�������'��?�Ё�A�}��uI{��<���b|A5�&Wt��l
���Z�s�T�wr�6:�0�a�G��^{u�r�0���i���EO!�u��r�<��v�2e�L�((n>;���{��:z����Y?��qeeu8a�3���S��c6F)W(J�O K�#���*VYm�W��#���eP�U�JҔ� X8F��8
צ�O�˸��ip{�������u�z�]�$�D0I<����B-�0I��1�HF���F{X����ܭ�#7���~Y�����\�%�l3���ȇ9�!��Bb�v�Q�B�㉻�|���&�:c}�Pt(�Y���H�خ�C�������
�9��|�D���ē,��K
I�v��:��\�A���9]{�16`^��(*V�8k��Ԏs�f'����e~���^�W�w¦���bk�W��ȩLG�7(lt9�s�}2W)�\�q)���{Rm]�2�9�����0(6)��c[�kR'�[�
�r<_>�S�]>�wy�,��s�|��F���@F��*=&�[��&�R���փ2!�ѻOpQ���cf�y�*�O<�D��΄A�%؟���}� 04k�>�h��^L������?��1Ǥ/�R��0���I�9gƮcj�K˭��E�t�G�	�zR���A@,���+
E�Z���ao���-�̧=	=��󌌜���j�9�ǿ�W�<Z�*�w�.Č��y@�Ff~"����#Սu�ؑ�i&���ï�Qt���G�L5$%����>�gpy}�Z_Y�^ kr&�c����'���J�Ub�bI�ҹ���Sݕ���{A�b���t�j��{��e�l���G��BRy��V��t�&���h��Fa��Br*��S>e?�'y�-Z�*� ��It{W�F��q�:ߕ�#Gq�c��WK6h��Xuh����	I��}ܼ��ƬO��9(�Y���Vt�`��Z�OMUe��M���"A�9�HA
��|��q����+.MY�Ua7)��I�E=y�Iɫ1��8&��d	��nu�Y�<�c:�s���B" �Ң�y:v�$�i\>E��WzUyFP�� �V�U[ 3��T�����}�=���V9�=)��
Ű�R�U��
luo ��#[w������$���\^��[Wu8o6��}p���c��C\}l���*{������"��
��^##�
�ԣ3��O8�3�<Z{/����7�3����Ð�#:�b�R=z,ƭ
{���L�I�u�7�ϔ�cD `S/e-3�5!�烐�k"��=��e�u�=>�He1��;]x�T�'�R�5�8Y���!%e��|#��F-ޒB�� _��=�h������yr���\<������*�u�a3"QXDz�{)�����R}���ק�e�䣮mb>��ҽ�|v����ɷ_�W�D�Su�|��N�� �0�0�57���AaG��r&t=��о�bΜ��,n���cv��".JL��v�� ���� ���?��q	��D�:����d��`�#,]t��a&%ٖ s2t��e'S��w
�t��x��ܑ�~3��j-�K��l�lLu�u����RN�bJ��I�d)�T�*g����-)kK���)D��֭jQ-X)V�?)F%i5:/�bl�1����:�d9�ٷ�C���WhE��Q;���ݪ�=q����#k~��ͫ��R�S�b�a�~5��5و7��I�0�0�;E�q�w�8X�D��7��'�|R��4����LX,�E�rKaZKoO�����]).���ܬ��0���d�iZ����E˘��}���ЋHo7N��}�ʦ�?y3�� \/��r�4�c�=�Hy�IS�L����/q����e%�\�=�1~��U�-:Bq��<��@��;��Ě{R�mTj�V�=�b2��L)SE^��B�ִj4��&����׿>��+��R��p��ʻub��/c`|#�Ŗ2-�x���K�]����������]U�6��G}�M��>�	2����)g�fuS��
�gu��u.>]!�C;N
�+p���+9E�?�8�t��v3e���:eQ�BU���GZ��Pu��9���Nu=?O��E�O=�TL�Mb%�5�+��s!d�Q\�<��|�	���b|'s�f��A��I�G�LC������{����SXtQI7g
��[�k�zT����WCĵK���-��vU*/������C=$�>�#)s��C���Q�8�O�3�T�E~Kqh>~���vb���n_��Yh�@��ԯ�*2�!�D`!����3�<3�|�����}ᛞ�
i�e�pN��ʻUM�G�J�z{.�j7�nW]8[���F��V����Zd�r#��A"��(���A�fH�D#1J�n�꿛�Pi�$BF���u�8u4��,�È8ыn+̘9�\0RS9�?Z��00��:�kr>���2e��e��	e�,h�/�
iv8��&r�R�g,�� �A"&z��K9W_9��0���,D���B;ҲGv�y{�t�[c�a�`ԓ��`�1-=����0c[,��NZ.�#e��T��9N����J� ���� ��-~57s�͂�B��mv4��>2ѤpH��e�]&�.:^����7� ߱8V2vH�|X�'����z�<�4]��rVV�@�RJ]B������D�F]�"/V�ǻ����5�\3�3kM�K�q�7�g(bdcY�g��
��}��r�,�)XP���曷�n;���V���DKE���v���:g��1�/�"9�	��d�D^-���!w�yg<df�d�{�u�]��2�^b�a�u���zD���Š��G~a*T�������e$��n��:o:�3���Es�� 7��ȷ�OS�ːbɰ�����\����U8�o=�a.��7���"�aey;0�;W�q���m�X�/��]�j\y�>��8BO"D��x���o��5��'< �"�g�,� GLY�_�dGW~�i����T8�R�m_1�D�sQ���"J�/��aغ?�v��b�-�n�˫�G<�A���n��,�tlC1�9O.$?ٴ�ݤ4`����w�\���X����6'ho�ꢀtu�[S5UxrV��(j$�Y��[6�pCYe�C
��lG<}��=�ܣC�%9`)�ej0��v6��YT�MI-�F.U�7b��϶�| ����d�L�{�]��Ȅ��EP�et�p���X�����;��.�������G��n��R��#�èֱ�(��PL�K*��[�b�%�詌��L=#W�v�(��+�jWK�P�
p{�}^�q����u��A/�Vg��ý�:>�����޻(���'��?������S�C\dm���>f�a."���O�n/?x�N��vς��<�{ǌ���AJ �F7�$kz5�A�Fi?)�|߅�']Am��x��D���xoT>dn�&ɬ|�7���Ê�w��/~��}h�h���0)��mn&�L�{C!k��{h(�U�}mH3O�E�)����/wL+��`γD� ��/�|����]�:�[\p�����/���~N�����P�fe�=O�f�.��"�uk���dTt~�Yg��q��&J�A�A���Z�Np�VS���:\��QmXD��kl� 6B��}��W�S��,�:���I�����t��&���^q�l�A��v��D�/~Щ,%�ck�=�\U������q����7G�t�_�Z�U8U���`�x�2�,�¹j�.�Ј�]���_|q�7c	�+{��^6�ʃJ����Mu6=��۫p�V{.�s�n��a+rf���R����UXD�\h���V�W����pҡ�i.�ꪫ�Yg��|\�z
�)	^�U�1��r�3������g�\05�.L�H*H�SO=�f�޲)ௗ^z)�Ӈ5�|�dJ��!�@������U:b$]����W_��#)c�:_WWV�X�[71�!;�b���#�+���y/���&��)h�z��h�j�Ê�]w�y�喫�r��snٔv���2�3��j4I�c㇬84�}����91g	{��ʩV&�b�)o�T�����E��w�|��^.OB|_�����cv�5�l��&V]�����6� R�%�Q�����o�i����d>��RqТ�"J;<������N9���ES�} ��/���GI킆~x8s=�lU�6)��]C���j�5�b�b����｣i*Z����I�c��s�SW�N?�p������{h�B��Eo�A�I?�� ��_}�1y��*L��fcH0��4���S�LP��o��u��	�s#&�T4�Cy,��-�A&�����}��&����(�M� p�`���Tj@6���׼f"��m^e�R��_���EԐp*�?�����-����o\�FW��]^�܄������Af��v��@<��/�r�#���_�Zx��q���_�8��g�yF[�cu���K�~��*�T<Y��5T!zv��7�6�Ua3���L��T(��n��i��s�.+���^	ޫsi�~D�[���p�	����sr�p��@s�s.�&��qs�1:Znc�C$�8�e�wVD9$$��IƏ�����)y
�SS�Q��;.��F�9���Ut�1 fh�������/�K�P#��7������_��=�a)��*'����~�6�l##d_Btpp�*8�RnȈ}Q�*W7�7�=��z�Y=Z�E\QxM��|���k�7���C| 4��~������Ҩ�Y5{n2���p{��S�h�ՓO>�k�E5�KLgHNq��7K}���G}��SO��O"rTUn�j7u�Q.�`X����qY��B5�#4d�t�K�'GO��}px�'����#�چG�Z�+q`H� u�t�ז&�b���R5�a+�?��f,��u�L����h�=��SJF�vgB�\���k�x@���������gU��35�Iᖘ:�a�Gq:P
9&iF:m���Z@"�JU��Ü��1���'�Mɦ�ڲGռ�u���U�T�����dsґ	�0$a�cz�������^�+�{�䍮EaЄ1�뮢I�w���� f5':�y�$4 ��_�KM� b^xᅘ���gC�8dqC�T�[���.�,4)��"�p{�*�=v
us��O�LY���E's]���� Z����B.�(P�DN�e��v��jer�'��o�;��N;��n�B��5A"0ج\��=��M���g���.�,������\��|>l�\�I*9��
d<�v�&�t��z�"B���ܭM*�t��G��`qJ$�M@GhO��zOo/��A��>�&�����DF��T���1��y�7�[�ƔEa)�o>�v�6�R�<��4uD�hs�O��}��|�P@��(�<9z6\n`��c��cgO��	U:���#�8����6	,�r��;�8PNO��G����?\e�UZh�Ժ�1���s��#�<Rp=Q�:O����W�ݞ�SCU��P��d�f�.S�=�r�-q-R��ń�A>B��9����N���S�,�ͪ���1�����-������ҪA=�L�,�ڎG{vjx�z���D=�hV(I&�_���}�݇v$�C*b�
!�k �ozӛ�hr^lv�E(�u�U�-e��ʏB��w��.���}�7����nĢ�vzx9W^���򓟬��ڛm��}�a(6��1W��G]�)�1M� �������r��9!�ziW$��Ą�?��O?��Oz+{s�n�H�����L`�����A���h�����?�S$>�@k3��O?��o{�e�Ym���٦Q�j��r�,0���w�i�P��9M
r��RK��U)u�dM=��|�����i�,B�4zؚ��@�����O9k����}�P��������"�D��+��� �#�s���O0��fT���<S}@ƙ�Fm��v�y��N������6P�p��P��R������������8��wn�����k����˔����	�x��J�T����d�NkT.�읃�Y)�i�Y>��s��c�v�~�O����u��ַ��n_q�S������$��Ö��Ԉ ܎��җ��=��V7���(E�@�QT�ӥ�^
����	�q���C�v%�G��\�Գ���$���|������K�AC�+3w�Sζ��(�M6�$����}^A��.C`~0},)p;�ݾ���X�0'H����'_4�n"��G�y�ӟ��vϼYQ���]�G\R}�D0c*u�a)�gv�o��n����E
�c�!�Ц��#�� �!|�{Y�C9d��V��"�D�`��i�K�����}�馛�ԋ-��
�t�� '
2*<sl���v5�t�UW���ރPe��?�Q����L�`\��,�ŷ�ŀ�u�]�;O��Sk��+�FX���o���?�w�Q/6��86B�c�a�b���-e���C/)tĻ��N�.��b����0�~N�f�M8��ͣ�]��>��
DXc�5 �v*�@>V��|�+���a��;�뮻��o@tׁ��ӎ8þ�����/�V�p�0�/������A�G4���=�|4����=C�X_Xt�p�W���W_}u��|!3r���u�j�s�9�O��ȿ}b��x��\r�%�_���4j�HC����w��u�Iu�z����Ex_��\�רΙ��9�,м`Q����/���f=+��:?)��
�*C"T$Qѹx�B����
���*T9�ɋ%4�U�0�a�=
���Z�z5қ=�����\�,��z�'(������W���O�S���4�n��k_�(/��1��p���������a�^jA��v�HM?��E�נHk��wWJ�C
z閉�����C��Fe
'y�[��H��9��=�:�\���^\vRo���禛n�c�]��]��ҵ�aJ�C�����:o7șEʎ��>���f���kR
H�P:��_�9B�awu�x"WRJ�_��L��O\�#�8B�4&)��%,�I1��_~�]w��'�6�[s�A�na/�䒸�IQ�4���2�5�\�A?�'�R�tȚ2G��g)�9�ꫯFI~�s�{�_(��P}�D"���8�V_��������u�Y�N��h]���-1a�,ݞ�]�:Tt4���׿����l�7n�V���,�H�W���; `W�ʼ�E�*V{��@:>򑏀���~׋1�{�|00z�p���6�WEfaՅ��e�ڶC��N�!?���B!���UTz�q!i�o<�_��"�ؒ��iYe�U�c���D�7:���O<��,�认|-fޱR?���^ziT��'x'�I/S�,4�]Ԏ�d(�e�j+�]v��я~c-ވt�pp��:�,h���{��I�	W�׾���U\$e�WtHi��|�O�T 4�Fm����[7��c�=M�瞩pζ�y._�5�u!4���S������!���3�� ]'Ǉ!/-:X��8o����&��J��<�`�!��=xk1�K�4�4.���H QT���%�����B��.>H�FQ��E��� h��\u+�4�:���K/��}�{J��S���"����y��be��6�8��\r�Ρe������v��"sZV���g���i��)��� ��_��g�wl	����Lx}�p<lC��`* �{p0r�x^��WE�j��b;� ���x
%_��/p�Q��g?ː6�l3�z��Ei��>�v�:5�����zD����SN��Q$_�ʪ����<��/���W����3�pc@��=�yxHzR\��͘���o����g�^�4ğ��ۋ�-nz'n��o~��SOr�±���x,�6+۳^��뮻�Ǯ��J��@��V0�B�u�9�9��CT��<�RN�s�.N��S�l�w�%�'�������P��*���k�Z�����j+זM�,��aMy>9���c>^�G����<�$��8�����Zu�� 0�	
���aV��3υo��p#�j���ܥ\2>`!�*r���]+e<��0'�AOh�������U�Q�y��G�J�Qu�B����_���+5��t�{�ƹ��릌	܎F6�=}{)�*C�}�c�o�y=���$_"�S��?7�ʅS��I'��+>��-��26d�\��$����O�s]Y�#�){��x�ް�"�8��n��hU$t"~1^1p-4�~����Ԝ��뮻X�.��εkl�{��Zw����vd�կ~�v��ғ�h�*ruWS s��~��᥶���⢋.BW�A�,�d���  >����^j��\�!v�]&r�1�0r���G\bq��������|��S@p�Psٝ+L�W��I�
 6;���a�q�[l��h�
�_�$�v����pg�wϪ��ǿ���/�Ä���*X���{�.U�<����~�4�TV ��z�;ޡK-�M�;�  �L�&����R~u�7|�@io��1}��V������>:6�97s���A.T��{��ַ�Ȉ��U�s4���n�f����P�!��/s�:��v[��:�߉�x衇u�Q( ���6�v4�駟��W�
~z׻���4�M��A��x rW�Pਫ)�-D��%���ʥ���;�3p*x��̅�-^��G;�-4�ߨ�T��U\�X�#�<�#/�͊3�m)�?��a�v��7�9�(ϝ�/�৞z�6U%����82��{��Vx��o�l���WG�E��\)�a�A��R�� 2`�,�{���r�pc_���UCyJQ�2=Ҕ5�����"� ;'u` Z���N��e�]��:�qA�A� <A%�h�]w���c�JxY �}�Ѭ���6���<�=�������۝�'K��@q��1b���1l!��U��'>�袋*�㠅�K�p�	(A^��:�:4�Ԅr��o{��`�;�%�xx�0��;�����d�@D��}�^ j�ueo��&\8 ��ˢ+�q�`E�u������GzvsAO
G�q����$�� ��D;0����2����V���䴓i��S �o|���w����0�_|�7{��WÍ�ܾ�r�91o�ϙ!V��=,W7��'�jM���瞋���>8��*)r�0wT�\�͔wB�]S�+x��CN�HHS����x��U
��Z�6��}�^��(�ŵ�E��|[�49�sXY$��-�Q|���_,�^{�;���;��t�a�/��&��OF�PR8=99u�mHM��ίXMG��Q�[�k;Qz*ԛ.�7*z���� ��k�Mu�a�"5{�8�@s�Q'�E
�`���Rz(�<����+��¿�eɒ&F�c�S���A>��實&#�Nh�����l�$o�j
�)�ՅdD�b3��ӡ/�ԛ��fT���sGd�?�#G��#��Z; `=�(m�馪�_�zA� f����6J8Ff������G>��EXu�U��#t��y;SCc�۬;�f��
 �CU���Y����Չ'�H��rK��*S��0�8c%�P/�Yrm(�f��3�*���PMI�E�v������+����4��3�<>����\�:� ���ט���-  %������梤�����i��Xh$���пh�L�|��z���A��?�裬<�?�Ag�ᒋv�F�0��~�(:B�]��?���ޣM��ٽ���\�DJ��k�����oj��ha��D{�m⶛������j��+�\}��_��W.��b;�G�\�44�T��ң�Rރ�W�e�뮻���Ք�G+�L��<�IC!�H"���Z�o>!l�ͨZ��7�ycHh�+��b�u֡�W\B�l�Vf�R�R���ͨ]ƞ@��^{��Z����x�`(�j�g���d���,p��0+���kw��Eڙ�8{�=+^Ktn!r��dr��L���3'�� h��6rJ�X AI^ʢ0l�] #nčmN�����a0�t��!���A��qi0!�l��4�~y���C�'�ÐK/�4o��=�܈�1~�J6���.=��5���/�jnд�V[MgC!��,)=�9	�kӹ��*�$���#�/��e�>t�V�!U��? �n�;����v� �j��йt#�!Ԝ��M���^L/���f�m�C�u����|çܤ�uf��̟��g��m�Y`�ӂ��9�9�܏����pXn�m�^RԖ����_M%��Y�nS���4V�x�+^��b�R��!���)	�$F�Q�0l�?��D�UVY�Za�qR��j+~���z�15e�26f��_��a3x�R�:�3�*�C`E�d��4*E*-5�JD�[l1ݍ����S Xr:�w�u��g6e����o17�l3����/�~�vzfR�$D�pŧm>�?;߁����g?C�#��xTE�XM��qD�|���By�H���G	#G0$�]j��C&���Z��w�M�s�c�����g�M�9B���R�|�a�g�G���hӟ�@�X�V�
O��D3�-ćs��g�d`3�����ޭ������H����iW���y:uNk��&N�p��.��ƈ1CpU>쩧�6ž�3H�o~���M��p;���FP%dG�4��~�7��?���;�<�>�ۇ�:���� ����uȗk�ʿ�Ǡ�S�~�� $�"��=>�=̇��͋�`$���Q$�N�T�({8��)�!��e��kg1�i�Yg���f��4���)���rq�.���6�3:��X-�4�!�T:;�BQƍ�Xг��0qؗ����K��m�\'�����-EE�`>x`���*X��If�9U���ِvTW#d���!�vh*'
눾 �j�`�����|]e��K��}����w��YDޢ��ű��ڟ�jYA�?�� 1�3e�iQ��I���H����R8��+�Δ��"v�Z�-�l'4��Pm��\n��~V��b2�V��M�Vʙ�4(��¦q���Ɗ&��2��Iaz�Fl����Ԛv�R��x�m
��B�.�\����~%���B����6�b~�=�X-l��憸z4/�neS�t����CL^�����h���|�zL���T�ҝzՂĄ��?�iv%�i�&�iG��J�g�v�l�����ȱ4�T�mA�v���ph"v�u<�YG?��c�O5l���DpEp����P]­�y�[!{�4�"��V�6ny�!�r��yhmj�g���p;0��SNq�R\���4��ݱ��_�8�/]�K��\��u�'�b�v�פ��\r��_!V�|�M�wg��'r*���u,p���i�C�f8+I7�kj��KK�8������ʀe�uĿ81�N��(�UQ-�A�N:�$��S�����L�Q�)��A�U�C@ƺʅ��䴽�ÜB�`Ӏ˺;<e��H��?+�"�%�6��	���@��~���Ga��G����m0z����������i�s��6�7�7 �]Q��Ue#1<>�&��|ϳ��a8����_���3̧�$�1MH�Vu837Uf'��B�U��n�O*ǔ�⭔}}I�A&�=rX�m}_�����"�P�V�@1�̣�lm�a�I�:N���D�4���!�iwBܭ���H^�z�9�
U����{�d*pn�p��T��i��N鬦�f��=swb,�7cxv:��$��BR�Î��s�Dw"�6N!�A3����͜faC�u����֭��N��gUV?:?N���z�u��*pW��S�11O R2�a@#�$}��XQʒ�b�j�GS�,&2�:�%=�V�d�f��|,����bqe��� ��� 1jѮ�vҔ��,:3�5�O̡�7�8ކ�6�ٟ�[lnd8��Wj_ϸ�~t�:�� �X�	�U.�;��:�N��ɨM5W��{R����|5�A�a(��O7�x���O�u*��l��a���[��g��O�{��&��6-�j5Z2�ݭ+�X�
z�Pʵ|͹��Ga*p�6}���z����{DQ���)eV404�	[dT�G=����:�.������y��w�Y�jJf��*$ť\�HJ�����о0p���!��ˤ�*�]��,R��-G&ѿ���=��L`��u�iTB�C8�[��-r����;T�w��u�PM_s�tr�	z��*������͝�I|���1b)�'�H!*O$e�����Z�^v~R�)S�aQ�ϰ��߉|���D�"��Y��5/�V2���j4r9;73ᴱ�v���22�����{�R4�|r
F���A���i[`�y���I�E%G�aK+xvu>�Y%���h��\�9�"�32�s��g��S�ח�}Ⱦ��[��s���R("E$W�����o�L�ǊC�{NW�d�_g����S�*�xUZ1��iq��{�g+èǼ�;G~K
��6gC��K�,�\�^@-Dj�n��h]z��)����S�U��P��.�a��T�*g]�4eV;�#R�g�G��b�K�f���n�T��́)���Yq���T���zH=�������%�#��j�l]�U8�~0[�o�svF���PT�����S�R�M���XgF��i�4�1�N��)�80kZkc�9���B�t�_:v"_�cy�[�EѬ���{��_#��;Vs�I�b�˸V�y;��I:�d�a��ɩ�[���D.A����ރ�=f��kw�:��\�b*_f)귚b,#?�	���:D�zTRO�v{Ҩ����Ls�
������ױ�D�\�h���|5�l���L�D$��i���.���>�Z���MZ1��aw�%ueT�/mP�ҤL�����J�B�=���O9|P<&I���y�J�0ֿ�^)U49~v�&�&�����Z���x Fl2�Y�ڦQ�î�s�_m�����Ӣ�ܿ�v8k�^�L�Tz�d�)b�4���c)̌-R��sڿ�5Rc����z���Dh����B�\c�)�d���֣{��ZQ����tM��A��M��hٌ����=$���j�N<N��0o��)�W����D1�h�����ںN���Jj���tu���6/k�iu�lV�4��#���k�
��Ϯ�7<Ӹ|�(�3� ]Oz�J��?�@^�+�m�kZ�ڈ���GB� r���Ե4�N�R��wt��9v����������ᴠ�U�EΪ��S�^�̀Y9���o�Ɗ��S��N9�S���0�K���v�mq��A� e^q��pg��z�N�͗�y��4�x�̈́���y1Rf�v�D��LZO���R��%)dqD�����D����M������B��\Lml'=K�DA��J�h��Љ&��QN]1��e1z:��y�Hd��[�iO�.>������d��~��֨�-pm���1W��i)oci���5��59]�Hq47�����|�������y��8�:�����"a���V,Ӛ����cm�,@�<����둛O�d�����S�c���c����z��g�c���vp$�ŵ��遞�/4֥�[�}����H�5�Ҩ��l��~tn���C<���q���ʞ��WkB/��)ԩ�N�vk7r���X=6��~4�v'"~J�-��_���2y�EW|"\�) �egi&}�C�>�Bx���(��!Q4Ü���d�%��R���������{Ē�t�BNzL�Y�D��E��k��^�*��3�#���A���p[�L�ma�\(��ʹ,n���a(=�O��	9�X����ު�Hy����yl?��ů�4��Y1x�촕C�UΡ4�W��� ��?��FOYD�6�%�V*vfcr|��w�)9�c�4D�_Q����~Q!Y������U�����7u/�T
X��x�rڥ���Ī�e�:��F�e0$��ȗR{A-��c�q�چ����boq�"��g��𐷉⤦�D_z,�͊�\����7��-�k+��Q'W�53R^�:D���N��!*��g�2��螼��l�[5]H>/R���G/�q�'�_�F�x4R>5����|��9����9��z,�y�ޚ�h^h��lE)�ı�A����We=K��{:ס�#G��X:e�l>�����a�^�P��GS2ȥ����5�����4z��Ra����i+6Z��O*��=u����-Q�ɱK�dN�L�����lR`����]���`�=�*�9`"O�0ӧ�����2z�~lZ9,�u���W0�-�Q���qi�E"�D��E�:�v��]�N���*����`X;F�CmG"SKi)�v�"8�5lO�����3�f�M;*��*bo�C���ss#˥,�=g*�wV@�u��8*�k%����|��0��z�ӔQ�M�т3�u���(��uU�9�V`� ����Nb�]�l�ZW� /��%Nf�^|�Q9���*z��޷���(EU㟧���������5R�2�Qj-q�"W�U���3�n�D֥0'��mq��9�XLV=���뇞�<ݵ��f�KT��-Z��3)Wuut��'� F0��ݢ�L����]QzE,��kQ6��KSPn�h`�p���ku]\���g����x1@d,��L�*�}�=�U�m��-Jխ�]����Z�m.=��b������4����>��U�{��_��
Ug"0�iA���fe�\j~��`��3	��i��&Z��%��H/y���"���P�kZH����jtg6�5U��s���˂���c,]*�8����hXW��Ǆ3B������{`:H��1��E���Y4O-nJ��W�IA����ÑYm�M|�j��ʅEw�1Fɨ�[�~t_�y�T�pW�(��콢�BS����O��$()Zܟ�Fgb�)g��E^��kW�2]�{Q�X�Ɏ�G⮊L��m0z"*zw&���A�wc��r[�����B�:u�S"���a!�Dr{RȒr~�>�ʭb�,��y�|ե�Q�#�QS�������͍~R�+��F���T�4M��2���7
���F�Jw�?e#�o9�+=f>I�;��k<#M���FO)�j<u���ͯ�a-gT�xU��O�Dx��qZ�_�{YD1�۷�6��s�G���|5zB,e�P�R/�L��\�U������a1\��Lv����Y��#Z0�;�6L2�E-mn��Ky3\c�����sfl����=�"����|Ǽ	b��oM^��K|�yE/=���jtG�321խ��~���*v�Ӧֆ>Z%��t!��.U�j�n�[�e"b�=Vg�=���|8���l�:1th��w
[mE��Xn��	?ck�V�F���t��Ě�\����mv.�/��g��%�ʊ����1g!���2{Y�!�ڈ�,(�ο*�z턚�*�6h
�[����bX|�w�yU��&��h�'B�>[h���Ϫ��˪F��o��j.#S�M'U��G�n)�Ζ��3�x����*��M��^���vn��LggE]c��ŠI,����+#�)�J K)�j�?�����3ǉ,�"�n�M!�����5�p��QW�z�¥z�H��xXӶ�}"_�(�6�+��-���5����6$u8�!K��N�#t0Ѷv"�,G��8��g������-�Q�������?�+ ږ�{���`R�5ƒU@��mV�r�=���W�?�OvM���*���W��̓S9�Wd���/�gG��4�������`�͇�=�y(�껪��!�k��ڙ��JՌ=�=�I�l5��M��Չ��H9�T ��Ժ]^��5;��/����dz�oy�-�"��-)8�|�o����DU�7S'�]�1ev��Y9�� e�mOS���ƈi��֚o��EX/�j��!Mژ'^�;��[�j�8��U(CW�J��z�� ��ؽ76M��x���W��2�W�*:�G=�+��G�$w�U��A��kq�j���󖬨ߺ:w���G)�֍���p���Rw���k�	���j=�
���Z�5�|�[��t�1��㕔у�OSe4U�zr�O�x���vk%`vZH�aqg5�A�z�4:4��6��|.7��~�������Wq�R#q�fKݴ��$�{��#�`��;��$���K��-0�>Ҧ��v?�=��mh�Q�\�������
�k���Q��p��a��#���i8~易��d��>v��lT<~��R��D�١���P���&�m�u> ��]����"�)����LAJF��=��\%��!i�G�ȏ�Ob/Ѧ.�#Z���7%g�&�t�R\�|��V���(V����L��MAlǺ�U�����-z���P�\ԓ����տ0�#�)�@�RȚ��lc�}��K顿�b�8�jT-[ l�O���E��&��,�P��:W!�%� h�S9���!���lS�4�����`H�i��ey=5	�<��eI�j�P�w���� ff�
��9-P=���"��ϓ����х�J��2�C�*��G�8h�%�e��]����O�]F�Rb)�nM�]$�y;���)cho)8f�F#����v����D�h+qk��M=��/e	2ޘ
�;.��~�͸T�R(Ӡ��>���)K�ō�a�����H������oU��m��ow���H��w/��M�?5�(�M���Zh�%�Xf�eX`��[ny�'{�'�|��H���̑~��/~�_��W��_������K.9�����������P[�iQ����
����|��[d�E ��{}�Q>�[��~��3 ŭS�(�I�/�8����>x���.�r��*g��}K�_���𒗼d�VXt�E��_�����@���9&��(4+�3�|�-���{饗�V?�0=��Oz��Ǉ��ZW?�x�2i"��d�����
����-��ȵ�3��Ta/Xӄ0	d�	�1�u�]�%��S9�;͠U!uޜ	n�9�ϲ�.���?���pl�3�̙Q�գ��1�������L�z��o��6x�����`Iц���W�-���L:�����?_qN�DI�3�Y	��t��b����*,1Ŀ��$M�i���hh_��u�)4��2�x衇P�<�4�c	������lE��]���|3�sR.�^r��x%�I�Q�b� 
(HQ�$I��3��$H村{������z�ջ��=�p�-��_�sv׮Z�³V�Z5y�d�ac-�}�OzV�ֺ�6>� �f�����ӟ�ĚBAO�v�9�%��H��[�z"G(ф�Q/p;�*r�O��8qݻ�l<)U�΁OXY��ˉ����B���q.ӫ{͵]��"�+��2���,+����p!�=�a��r=S��`H��(7�9��{�j ���sƦ=+N�d�%�D���?�j<��C�F�\xE�11����T6���ax�ð�?��J�;�/�`��B
O��tN'�a� ��:l�13��5�4��%(c{G�p;�V��w��4��;!�/�f)�&>h�0<|(�.�*F��c(��	���B+�l�-���Ҭ
��#j�c���D������!>t�,P���&{$�i�O�J��v(�yYSF��Bh00TB�9,[���CN�N�����,+�`��ovBA�vc�V�C��/��R��(1f��/s��y#�a_owh��g�_f�e 8��3���#��?Ki���OUk
�ii��'z2l8d��1�L b�a4������K8��ۥ�aB��!�aZw�A/X<�UYa���z��6��័Xn=����^p�W^y�D�a���Тg�io���l��ԩSs�^0�?�x�]v�?��õ���5H�@���G?�Q֏��vE�c�A�/������c�=��4��$ā��b�}�C�Z�,]Ί�t�M��aĸ�,��g�������;��z�G�j��g�s��]}�՗_~�=�ܣ��c��-�� t�t�M��+��	��vHF��/��b�U�Y+r�Dܢ]v�e?��C L��{��Q�O���K/��7�x�k�ꪫ~�j�a���ѧ�ɵ�^�����n�&3Mkhb��VZ�����k�s2V6UW���_��Ww�u�N_��^S�ED�]w�u��f�UVY��hva����|�͗\r	+kܟ��Vo҈�0��[n���Ù�����4G�~�ߠ˲~�q`S���dʔ)[m��D�2ز��)4�s��B���1(EWa�5��~��7�pC��8#���g�}64���-����e��u�V[m5�im��9�@H�9�'�|�t��>�M<ƏV\k��v�a�9ܮx�.�Ge�w�y7�x#�*-��ǥ���KCA<Q\h `72�U��r�-0��w��,�!��!~7@�G��9`P�%���Y�J���*��뇌�X�:@m�}��v���cV��e�H����Ha/»���W�����gF.L���sz����yj�
��qR�;aȍ���2�]T��3xȎ�^u�U
xy�_N�qRY�]g�uPbm�����g�G�����n��������OQ�V�֑Η[n9���g�|�v֑���OpBfs�
��۶�n;����ч������5���|����.�)��|�����W\q�ǳ�q㢡�_Cċ`H�S%�'���c�>2ˌ�kQ!nG J��aUL��B�;�U*u��L�_伣���few�yg /�ۥ!e8 V����Ũ�i��6x �FR�/Kp�}�1l2�puL�KCN$����Q�/��D�������~���vч)1��ńi 0��Qs��?|�nl`At&3W�N])��G�Q/�_t�t{���O��]t�#����~:�p�[+>y���wߝ���;�&^.��g��@�+�Cu݁�nC�R�7�X*�{衇b!4d���R���Ј%<�c@͎�C''m��>����3�a�)W������A#:?���:�,փ_*�fX��=k��O}
��_������I�P�(��?��`�LI$kz��W�[[�R�C�	���%����g
��]p�'ā��ί����TI/2������o~$'=��/�6�������{H1i�V�m�^��q����]��v$BO+\M~``|�':UH^�3����&@�#�8�5��o
{�ZzF���taA�>Aym��'�t�)�����X��I>a�C9�레r�-`�5���#�ԖT�ݲ����t7����/��>p��꬈��*3G����ߧ��a|��:2-��!<��&��|�Q�8��P��x�)Ad�� K~��p{�{_)�B���G��~���D��k���`����g�I�i9U0$��~�d�MD��H�5��۩��
�@�i�T'^@��9�;�	���y���K]�gq>��׾�5�*[���ʜ3):�,��Xg�څ0?x�)���\��k��`B�m��[�`B�����?�1*�y���)/Ձ��]0��1�\0Wai�
�����~���Pg�b���p���oE����d�y ���;~�;ߑ��m�{�� ������!c��8����"n��{�0h�d$�eiK�|������??�FD�����E����җ����J+d�*����	�����E�Ԏo���uI\��K�����'3FL�:��)��uPl��X�,M���_�*H �^Y�&ū�ךk��r��{�Ƅ�G��!J���fT�!M������'?`���� ��\f��9՞~�>�2O!��O����y�hfa5>�[$��A|̽p����2��,B"��GZKִ�קL��`lp`|;��>	0	����>��m]��J~��DL��H��)��s����j���2�3����y4��{��;�K�{��Q;����>n��~U�	�o�|�1g�p��R3�}6��`�n�AI���9�NȤ��W_����Zy啅��'I'n�4�6m�x���ː�޿��!�]?��Ob���|�NN)<	�Z!8P��Nõh��r�,��>K������N s�������.R
Ȇ/��/��°��\�A�t饗��A��JYE�9�Y{�5l�H�@��H�#	�����ZE�<�2g"�,� ���o�Պ�vue�]wE�a��\�H�|Y>���u�@m��t����1�eά/Ի�U�� ���N[�����L���O���QX摐�6�;�1o��p؃q�X}Է N�+����L��c>���o�x�t���a�pƃlHng�Zʬت�O1f��p�:��4+Dç?�iX�jk�ϰ
�: ����4�#�z>~� 2��>x��J)U);�| �|�[��ude�3��Hs8UE�^^ds�p�v�������7 [�r����}�c�WXNL����S�9 �f�}�e	 d�=�X�k��"��`,+��7!^����-�
�+�3��qא����v��砣�Z�N���/�<������r'�ք4����$�7P/ �T���ʀ�ȥ���?���=��1��q��.��	��f'櫕��*x���Op���kn2��F=y�����S�����ox �.�^�
��1��ئ
[��e>�C'r�Q��-u�Yg�����v��������7qG=l���7����%� l`?E8�$t��a�P50[ru�ǔ@�iYt���#���h�H��'ˊ��i(s�c�)��!BBQAp�k��֐ ��#�K�]a�
��,Ę�
��x�@[ �ֱ9!G�}�-�dH�Bl��x�����~�=�虑�������g����P�:;��n�ݢl�� �'�|r$��K97a�̫�����J9��FādV��j�4D"]�w�ygV���H�}
�WCy~�p�	��6��б�$�ˊםC�c�	  �~/��R�O��������	U�2�b����Նu��\�}G�J0�c}�
�Z�1xz���PA@e��7)�"T=:�7@2�1�l�br�	M�8��ݐhP�z��9��L����2���(7/$Ӝ���uNA�p;|�8�j\��#T."��w���?��vA�9͢戔�
� �~�V��\ʧ�?��k/>��(�V���_����(��"}�;)�@�
�P����P�5kg��_[l1dl�V��s`10��i]�� 4r~���;14՟�6��
�ts��Z��jE�K�HP[�ʷ�V��<��A�F�s�ֻl����Kx̝|�,j��\j]䒇#����vv�|�+`~�=�X`�5�\S����\k��+baVϨ譌�dA~�Z� "|b+��Ǒ\��YȨl4\y�R�yJ��13S�D���r7��a�o��00�]��,�X;V��p�������H���^!*j�BFZt%���E�;740�	u�
��Ede�U����I'M��Ja>���'�2��_w�u���A�I��ȕ�Գ8G������H�!Z3B�A�
u6Q��&J^Al0r�8�S�mO\�#h���p�5����|hUS��(Y\�+����Ɵ5��ꪫ��0?6�P�5=�V>��Zk�����'ϼ#�R>3Z���L���4�6mB�`�+��[�J�Q���m���j����,a���o�=������
G�GC�E� ��]�O���RQ$1����|��>��	���P�^1��?�n�ݹ���cs�5++�>=�v��,�������1�����%`e��?=�M���e&��cn���(wr��ǣ�>���,A���j4fG=�@O�7޸��:��W��Р��%��y�����<�\c�5н��?^+7W�3�.�	�`��H>�*�h;"�Z ��^Z9_�����\<j�M7��l�\ê6�2'O2f(ɋ��=oeU��qbv�}w�r1IU�/ib �1d��?���l�1���T`�_{�\��A4��_�~����sH)��)�/ݎ�T��z�e�$s�q����&W͊���F�/@2x`+��I͓�vDRs�1o�"u����^ G�ɇ?�a���w�2ւ���u�Wh�|��{q�T��)S�/d�cVO�&�¸����n�=����ܳ�[��;��(%qo-o�����K�e�]`B������D42��4�Z'W+Րy|}�u��|�J2�ܮ��s�9��=��vs��M6ل��q�a�͵�p�`��n���������9m͹zz�r�-��]����� xE��E9<�Tf��v�Y:ա��g��'��\�ҝkNK���Ƀ>x��7Ǫs.���yFE"]S�NE�:������ 
@�+r�"���2&<����a�r�����<�H)>�y��y:����ɓYMe��\�%�gl��o��ꫯnp��2E�h��VB,Y���H�T��N;�������׎�M��$<��[�!G`��,�h7l�=�����J���8E�����Rq��zȈ�?���g	?�m7_�p;��OA����B �N<�ĆxZYx n��i�E��:��cx �M7ݔ�e�a��{��v����̌�c���O?�t
Ĥ`�*84�sb���)� ��?��n�:0�uo��#h-�]A����!��R����;/���x-|���Wf�o�j��T�F��Q����o_���P(6�|a���_W����gLQ�^�?ᮻ���ʜ�Cts��\f�e�nuB�غ9�[ 3q����'_}�UG^Z�>��ϡ�,�<ZMhh'�����V�pQ�,��<
�e�P[n-��Ԭ�7��L@�n�l�ͼ���UnT���;�S�~�����t��6�i��_~yh͝��a��7���'��;�J��6�l�V<묳�����0 ZL���+_���)=�mXTӭ����_��!?U˴���d��;7��2ʐn����}�Q��?���)ށ7%g�����`�ظRP��g���D�x� k
���Q��џ�n�!dv+g��v�CS��x��@�[�zSR���X#x����+M�����$��x�c���Rm�A�C9���?�1eُ<�acL��RK-�l�R�4<�#tl�(���k����8Z���J'+C�y�4��Eq�ݦYԼ�*_��[|���b�Vu`2I``k\��/�\���#���1���B-T�M���auA\,��C��5�p饗FAx�&��>�D�L�0��W�0�o�5�l��Q&V�aC5\z�t^���-�q�aS��2�`5�s�98o��w���i����:bxd�����a��Q(���v7���+:�f��7��0L奰�%�u�Ӯ�C����z�!���)���n�Ī�\$�6�|����^{m�󵀮��H��:o�����sύp�����_�PR��K7��G�Pi�Td]�D{���zYxo'ҟ��=jk[Q�W0���;�.��WjsD��[o=)������]4y饗���>�bҤI)����M�\r�%��������2��k�#�p�?�䓎:6�'0��q���
�����	Go@pl�=
/�5�N�&�:�~#��ruE�Тh�[n�E�����/>��ލ6�h��W�S�vT9<���/��˥�͕�@;k$��V���߆ƴ]w�uQ�gV��o��2r��I%�z[Î���Χ�������ة��X�a�:z�l�#3�L	�!~+_�g@C�	n�1m�s
)4{�%� ���o��f����@��S��ho�����c���O;�4�ѹ2ԕ�!����� � F/zQɳ�n��J\1��-<|� ����p����W�~�.����t�CI�p�ҀBH��X��+��,�5H�.H�r$��,�
�:�k��@lR��:��駟v��9W#�H4�z�p�R&��9Ux�t�g�����8�O{�X��ZH�13C�vm�οj��V2rѡ	܅h>��I��'4��?�r���4F�S�N���k>a������[���?W�b�`4���*�Ԇs�k�ȗ_!������f�1_���^�䕳�>{�զ�XEQ�������+�� e����W\_��\E~�ls0��{��6G}�;�2������e 0���qZ��E�Xf�J��H\��-z7eį+��2�w��g�G�2 ��O���]9�[�<�u��$��ӿ�w�?���V�ư�E'S���G����̮~R;��-)2dx��6�*��Hy�����6�R"Mt����[�#1��X��,� ���O��|e�0���� ���o����:��������|�>�����W����g?S�S��k��[`تO�Z��_o��.����S!`�[�p:�I�r���"+q��C��a��AhL����ϻ����j3�3���j���3: :J���S[2�wT����I�	��ቇ���"��x��j�c�9�}�.a\+`A�_JG���l����jp���T��m��:��o��4,_5LQ�g�s0��
ɬ<�f�(�p2���_���Uq�"E��Y�Oa϶��EH���z��X
[vV�p �U�����y��*8%=�-�ۋ����5$�3�.F�F�UPW�!a�~,�\��n��eN�ձ�}�Cg�uVw�E�����X�}���ywpG��zȠ�*�Ȼ�s�=7��J�7�����r�-~�ꪫZ�������3�<�H��ދ�vƑ ���*��f�!�� ����2��j��H�Veڴi'�|2��²��]��:*��Fr�P�
xC��y��k�V�~H��{s�I'��1��P�K��E��@n��	�=���z<r��o�-�l�n>�]���|/S?���*�SJ �}�9�(fd4b5�*t����B��3�+�j
0�ȣ�>:,��`��i��XZ����)��W_x��g
���͗�!��R��O���{��Ile�|0��:�,�)D���b��I��Þg+���RcS�G�-}�
+��|���L�d�-i�q����A�����Լ)M�`K������a�)����Gq~+T)I�����&�$&�E�l��z�s�9'F����hy�>p��F���8A�u�Y��N{��7S� ��Á�Zpl�d�R�#JH�����Ϸ{k8�"f_i!�pǖ-��~�5b��BT����\�[�	���ڽ)αGz��t���)�K3%�"JݙU�h�L0i|@ޑ}~�0S�k�R��:ޭ]�-��=l�xY���V��u��-���,
�G���D�T���(��@;�2$��8-h|-�'O�0X����Aظ�ӰQ.ň����}��`8�%��Z3�UV̻�����Ԕ)Sn��&/q3����2�,#��4|K��&�1 ��#L���h���j��0<��U/~Â��qR�U!�5��|�a���p�@�DӨʼ����O��V͍4HBݬ��`�M7���/�e�-J�҄!!�7���va�Ѫ����9F��XX��XR�� �����a��b\�^$�>C:������J�ȎbQm�Ѥ^� �5d�-(dA��V��Bu�+sD��Q��m$WsO�0��S�^q��裢�*Θ�n�0�ws�>� �`e��.j.�s��RM�68)��/��R���3��8~+_")�c2�u�gԌc�Q��SO=5ek%iꆛ�YX��l� �Q|K��6
��[oM��P���nU����O���[�E8 ��h���|	����n�P���~W7_ޜ*���~0��-h�G���\�_2�����oC��Wz1>ݐR�:}5��������--q��{���5�(E�l+�`n�喁��Zj٘(_��>T��0��k��oN�H!���c$��1Y�o�&�f�W�����rH�R�s���<�|���(�FRQ���Eؙ�?q�F�&/�^��f�����n����ZeN��0��)�7�CԺ�"L���7,J�C���s���<5^�]w0>�]��KXheF�P���~?�|���RcMA"�3L[�s���jmE�|���1ר�Y�|�_�P��e�X�ai9����Y�3l�p���@[^TYb�v���a��x��'JK�Vaux�������U�Gs���'[��qF�~�4黓&Mrnd�/�6_X]���[ŲL�c�EE��1 �O:!�#��!.��N�_��vN�-�,^���{�>m+/o�T(��} �y����۵_�(1t{C�"�13E�۹�Qm^2s~��f}�Ȇػa����h�LPs�Ȩ��qHʓO>9�a�_��=�f{W�%�Vڷ�z+��6�0 ^��v�N���'��X�Ђ3SӀ"R��"	6~�UXf�I��˥��U�Rc3WÐ���gN�)�n��~��𨁊7�M�Tq;�weEԬ*5M\)�L�����
�P�0��b�����[!��N�� ���߀�5�#��O��U�e�M������Ji�?BG���v1�o��/�v���K����;�4���e��P�Mr��.�����ĵ�w+&��*�}�re�a�#����#�\��)�J���A�vri�v�no��E t��rfo���H�>ÏA�b��LY�袜n. ���ᔭ��@T|��.��c���Y��U5X�ۛ�Wk��BD0^h�t���i��e8�XTYg�.��|7�N��$_q��M���@�VD?����IL����s$us��v(s^�D/��G����_je=��l��I����M!n7�Jg5@���gwf	�&���hp`5��=��M��)t���L٪�.z�k�R��a
\gC5�*Kq+��'�!jk1<����hz�-�Gi�(~kXTMį=֠�Fra~"�s�y���*4�'�D�(B7�us���9=ײR8�Q�����U�[%��>��ɱ���oё�t�z)X�����I̔�ݹ�6�>�V>q�[�wS.�fC<�i�,���f���ض�0)g������%K�$dKİo��P�B�Ј��CPֆ��޴SR�q���`��}�L
�~B�̺t�N���\��$q�`�H�p-N����K�X�v炖yLS�y퍩O��������\(�Z���W�c ��	�h�Sۏ��C4iQ����l�����0�7?g
�M+A�guVF��\�QwǪ���#zy�~zu˯=�v>�S� '�q]F�A���"��t�ܰ�yR'��6�^~-[����z�j��1f{�3E�9�9�"aGK��vr�t�|�
]$R�����]��Q+�HY��@R��U��vH�V���P�����L��ŋ��n�i�|��x����v �5���g���5a���bcu%;��6Ǌ�xWD�d)s.���0V���uq������ e����q�cؔ#kS�֘7�N���КM��f_�4T<�^5�l~6{w�<�k�F���,�`�)��m7��� #�ڏzp!��e��Y4Ԏ���&Y�R	����h�fV�&>1X���L���s��f�[�*�����H!?�j�<l�p�	�R���:wyx��{e
�a�_�}3��%�:�񥴍6B�|0����~�{H��7�2~`R��ny���@�N���I�Xi���%McQ)�ޮ��5<��r���9S<��ʼ-0Z]�ij<ޗf����,���k�56u+��8t�v�
_�b]u��}X�D���B"iH�D�%V��*щ��n�<�g��$)���dc�8�nu/xL���[���dD��|��zЂ2)��a���\o���; �e�����h���)[) (������	����v��������.�a����E��r����/�N��2����gE�,jr���?/oZ���F�~����TW�yV>�����3�<�V=���"�0��^�~��%ކ#F-����`�9=��k����b�A��J��;eN��=���t>�=����d}�|�O�*�gj��)�ضm�7�Y���Ų��lG[!�NJG�n�j$����x�|��'����Mʇ����pH#K���^S��SOAs<��(3~�{�>z��'��~�)C	->3^��k�J�yz�x˘	��>��h�������ȄqH�b��,@��SݐL����+ ���Q�cN�ڦJU���=���F"eOL�_�k9������,�W�ӟ�^�����h�kz6�G~�q$ߍG}l'R��L-:��bE�<�Syq��g�}V[(N��'�Z�iE��� �q�T�_"&J+�t"@�'*7&O���+�!�(AqÄn{�1M+�5�b*a���������ԫ'S6�$���-b��9i-}
������)�,_Qq�n��T�@y]ͥq�)D1b6�D�U+sjo
q.-ӛo����5�\L,�a�����f��a�tǜI=��� �he[���Q�ێ2�D�x≁м�Qh2�7h�n6�z�/�sV���3.��ո���f�n��E++��B���6|B�s�9���h>��v +"����MC�I��0M%�h�&{�F���p��}`Ϛ;�暪���Û�x��v'�E��$�vq��3�"�nؿr؅/�!�&̐�V��7�|)3a�i�E���i��)ڏV�_��e"D|5n>�S�_+���j� �\9CwF�^�_���w03�\����$� �Ojv��ڲz�t�nvFTH�vN7���+�E�s���/�j�����!�/���o�Nv�F�w��x=x�M7�|iy۹{�J��R��9�\)�!1���auJ����S�%�wHX�\���8<Fqi��9G�/��F��XS��
�^<x�[n��315wST��p�pyܠ��ZD��o��O,X�APר�(��{�6m��לgQt�рF��}��ǂ:,gRX��W�d饗v�];!�*�$:-B-�s!��[Ié7%̨-���O��Ŭ���0bB��]%V�7~��>74TW(J������V��o$�"��r�?y������)� ��X�x@#,rI�ԋ{��K�����5�c�]6�P�U�[�2굒�}�TW�BL~��e]��hC)*��M��p��3=T���xڙQ5��	�{�6ݜ9�
�j�
����a5I4�(��=�����b�"��E��C='L�׻v{+{�	�E��2ˤ�����C��&ѓt�T��>��2����'}��4��?�<{%��,�$ǥ�Q��Sa�uh��d�-ݝ��)`/�'=f�o�-�d)�;\z:O�O�Σ���ɜ�Q5f�ͷ�/�9}�风��j+hU����g������ʢ�-�E8�$�ô�]�ΰI9{�..MW�2�o�QN�W�r*�������.jPR� V�qA�|6+)7�i���1�sh)��)��VޔI[bΐ����/��:l�qB�-�pH4eL�c7�|�����Ʌ� ,��g��!T���e�jBb�ãx��Mâ7��~SI�urF��&>��n���q���7�Fx�m�y�О�h�'��U�Z9�(�1}h��?���y�����q�e D
���~uY��eG0�:���%�V;`����.��b�5��JY�ᠭJ�U��h.g!��3ow�6�®�uo�:^��6�=�\��;�l�w޹뮻�����=e�T��N>�B�a�Z}E�X��S�L�Hbn�C)D���x���<�r �Ԯ��E�(}U�Z�B�D���#���|EMX���+��c�N^�I1!T~�yPe�V��7j>�u�]�=��F��򾒣e��!���
$9�����k���'>�8��Kk�8��[� ��V�)bu�ԩSS�t�S���y�[PU�JF�	96����AP��o����ET�����^�	bGR6N)�	xʷ�z+c�&��I&e�6!�lH���< �S?f�\�����l�A��k)�m�1ş�h��B�H�Sq�7���<H.���|�J�X���RiMvW/Zj��ԕ�p+���l���S��Gqۘ�2`�m���{ݍhS���7&���w�C[�^�ԷĢ0 ��g�}�x��6�a��	cH>�{ֻ�+{�u׭��Zo�*8����5�?+�sNkx"�
/��2}:�՗SC,�"�*D(j	��+�m���,F�j��yK�;�๠%��>�!�?�Cq��yk����AL&d�������9iҤ"T͋�-#���h��V	�du�����_�s�׮���类"��[��+k�[U7��c�":H�:V�!u	��-W�h�T� ��n�d�/��>[��)O���3�D��.�
�+g#� ���E���l�7�xu������}Ţڵf^�&mØUm&��vZ�Јۼ�Ϋ��a\k�2�x���|�#iH�ܡ^�&��s2�vQ���P4��w������?�`���f��=*{���N�u
�ŒG�2�q[n��t�N.��ώ92�%f�S;KN�ӌMog�0뭷�X���9OKZ�1f'�+DR,/�[�R8eT��nN��yI����ͨ�e�k�������R/�հ����v��6��t�Mߕ/�~1 e�Q��ޱj)����y}���N;�T��W��jN���ju�.�$=6��&z���<yr���S.S;���4�N!����:��M7ݴ�[�9���H!�Ԫ���?��>��s�{n��Hï`Q�\r������0� ���yב���|�b��g�i�5����l������	�]ݸC�5ǜ|��H	��l�9q!����'?���~�,IG%���Vkm��_��Wâ�E�������sO9-�F�b�=X9���&>4�% ��.���|@R��P��N�`�[e�����s�z�v�4$�`C˅"��
1l`0��hK4�d��:��~��t�A�_KF.�T��������Ȱ�F�Q�l(��n��6�l�R��b�$г��\0,�dU�w��_c{D4��
QIc֑ a��N;��W_m`r;ܩi&}�Ţ�.���|W�="�Z�u%�-�k;�WVSc��:�,4����S��v� ���DG�=,f��|�)�E/ F��cA5�������상��vNѻ�/���M�F�ɷ��}9��f�^|����Z������mta�y�O�Q�S�S��5e���~�N?��#�<�a��SH���w�H���qu:�j�����R� ҡ�F��"1�4��Z\t�E`�2�Z3@wx�7B��j����.-P�i9:��T4 0b�|�D
�@*���k���ۯ����9�Io�w�y����)�uS�����ӟ���j�|�`$�:�$���XN>D̢�`ߥ�^���z��E�~��D���x㍳���l�G�D�3EE�UW]�_�ݼ�ҭjn������O?�5�B3�+�}�I'M�:U�s2�1���
��9�y�J��D%HM|a�a+s^�u2�J ����r���tx���C���__�%�2 �K�������ۣ�,��{!8�e��j�j�)�"��qm��b��8��KYU��f˰��B|l�;� ��ɱ(�O���!.Bi��rC�������vf�B՚2\�c��t��/b�u.��{�*6�.T��aKǦ��b�}�z^p��w���r��SȀ�cػu�YG,�j���S�h�w�v���tɤ*H�F��:Q�,9�#�J�I���SOE�K=F�[�3!�E����=��n�b)s�\���aLk�b)n���;CN�G�J�b�<mC5�	�t�v��:�����O�(O���dШv�j���+����r�-���;������)%��ÎP�U�_S��5C���iW^y%��c��6��� ����F�7�x*����S���$NŚk���r��R���D�N����/�/Jr�J��}����=JeH-MyM�%F�&pl'4�����N�%�~�v��f�2 �ߤ�� 5*��6пbcq��>�V-s�)� �k��F����Lp��j�x�;���	'����H�h�2�]�5�=�X4���ϯ��`����_�d*���b��Wk(ˀY�w�qLx衇�N;��Җ%@Eb���E�i?>�����?<�C�w��p�N4	�,z>�<���6R�v�j� �
�w�m7G:S���"E��oў��~{�6�r��'ke'O���Zk���j��E�A*?����V�Yg�F�7��|����.�-��PK[���`���Na��ʜ��z������߿��b��Sp���܎v6 h�&�i���V;�b��ϻ�ah��|�_�]ф'ƤI��^zi�K�y��3�;�<�ȉ'�(���\�P�O�����?�җ������՜!JW^x��fk�n����)2���#��1TE�4���$�2�G;u����cQ�$ t��5���?�Z[
b9�U�{����X7��ʚ����(�����]��*��b����>�8�ՠH�x����ӆ�����?yn?�裑�[K�3wXJ�J?{衇�>�l��"l`vsb��	=�8��5����ɝ��ɰ/���Y���
B���c�d�M���ގ<`���Љ����,���|V�O��7'����!�x�	,5�l�����|�&��׾�5���Ve�Ws�h���Ot;0eF�����Af?�����o�3�<�c�N�-W?�>$<|�Wt�-];�L�}�uׁd$>� `|X�"u���l����N�P���ګ��z� �*�	�KHks�|����a'��0�ݎǲ�K,����uL!fvxۍ�U��V�e�Ib�	d�p�.Zy�B�5�l�b"�nkה�2AQ���I`̖[n)�d�<�JA 呢4��[�`k��d5a����h[�j�6���=�dɤ�M�&��|�+ȑ�P$c�s�A��}꬟Uf�o��2GE����<$'���G�z�q �p���`9����Y9�'�2��s���zN�4x��yRR���-i����(EsX���:
T�����P��� !�<#SԀ�%H\p��{��S��8=xm����3,���0z��a�'��H��C�<���)<C����z)����O~�S+��v�M���m`�)Mkv)��P���o~���^t�E�ī���@��������+z見����~�<��Sa�]v�&�Kwr���/~T��_�ZE��������D����S��l��@EN�вJ(I =�9A�X/��Y�\��/��y���B�L
��7a	��[�v`�b�
ˉ�/���a�c�9�s����s���e���Y����w��S�K��.�Q=�)�e�phբZT�%��{/��SO�X��&f{��WYY��m��V�M�W�������U�+�G{��������m�Q
�^�Xr��u�?�<ɂ
�{�յ��ls�%��>��O��t"�yz>�P��94A�����Dv/�5>BMx�8Ҏ$yGs��'(���ػa��xO����"�,�뮻J����/��:��T%#�Mv��1�4~�{߃�g��֚�w��U��+�����f�0Rv;�:ޔ�?�7��o`A�L�����H(xj:ু毺�ԛq���=pǕ��:Qʞ��]���@���;�#�PVb�\�Q��kF2��O�6-���s廽)�c�.Bbw�!�cy�
_7��&�:�X~X�EO�B���&���Yͯ~���@�T��C�a����>���U���Ӣ�P��������\�̩ݜY���;�S��=������b�_��W��g>�9�3�sY�h)��
�����l�q�>�n���N�Pe��cXmq� A+���y��nC�"z��-eua=%n�]�j;LS�����\t�E���~��B2~��^<^�O� �B��kA��ѪD+���o��Ƭ��!I��|��"�,(..<9��W|�F<c�x@�
g� J"�k��v�	'�cc6G+�0�XQb��ɻr��v.�����b!�>�1܈�jM���H4&&T�N�K�Q<C��(y�0���,���(��t�q��Ͻ��{����F����W�ڰx�����?��{��~)5��Bi��~Gy$����m�2�:p|\դ^��0��#��9�	�š�:y��V�nK����qZ4��D��U����w�<,F��o)lJ�P��k�Ac>��>/�8e>to���"3x,�XL�2Yg�%ۭu�n�3p����GB�����=����/N�ꫯ��m|�&<��U&n��0�])��W��]n��F�5m5HW�T�&xw0�}F�g�套^��}���93�pI�HJ�g5u.�	��-�l�:���2HVV�F�g))/+� K`t
٫��xE����瞏~��P���v��.|��c 7���hν%�}@��\rIo�X������hԖ����Yg��W�v�J\��F�E>��8o��f<0���K� HU䉯0�v�I�טiœ" |��5������@��}�_<����kR��먙ڏ~�#�@�eg4�!K!5�Q@�e0����.�ձ��|��o�Cx�G,�R�+ǘ�ð�9_2SyG�̅���r��4~�a!�TE��z�-&�!\X/\�x�X���-��g�ceަW|]��ƽ}�9��1>(���b���A:ގ��k��Y'WT�?�S�������ە�##*5�w̈�<�@`�6�9O�����E�V�[����/�1��G�V9�p �ΧL�2�V��
����ƿ����H;'6N��0#p*N�&An�"��w܁z�o\i����h����bL�O:�$�a.��p���
,����������R(��*�l��w�y'��d�N��"��lUM-��(�b7�M���h��?��]�*l�\!:Un��x���w]���O|�M7}��_Vݶ�n�5�c�*�j�=����o�9s��</`��O?_]�4p�w�y����0����s��(�c{!g�K�_j ����+��B��S
����g���Ϡ.>��O�����9#l=��ApE��L����������zx!�4i�o)Qk�4�Ĳ�3H��G�oqʅd4*q;��C\-�������`��� ��kB�K����N�x��
� 1����� t��h0�wXVެ��6Qb�VU��D�l��믿>�P��A�T�%AZڬabQ�k�#c#��݂_o���M6�d�5�PD��ӯ�k|_����<-��� `~�a,�V[m�*"�NP�8L�9�Xqx@G�:�ӶZ9O��OF;l���뮻.N�""�-膞���d�����B �Mw�`8&��\m���I�%G�k��[n�jc��;Ĉ�{;�(G���?X,��~��;��K,�PY!y#��J�t���A��R�%Ph�h����L͂��'G��nGB�n�%�||��E4&����F�ֽT�
D�OH8f�����q:��c��*[q�]wA���^[��
�p�i�=�\X?A^\|F��B�-v��ڱ�@Ft����nU���xc{L�F���S��k�p�n���[0li)}���bB.��"<�wṙ�D�p��Q�ʷ�n;h�wa��M��\r�%Jz�6��IH�g�����*�%2�UM4����f�gB�[s);r�D;C�����B)�S��0$D�&��w;�m[��Ո	N24�'�����0��e�*� ������!;E�MCjS1~���ᇣ�M��Cw)�'!E`YD:���+u�'���P"i�������(@^��z�!uE��Y&(�L]x���g	��b�o?4T0C@�^P �O�2�+r����WDC^w�uJ�+�YC3�y��t�$���k���12�E]T���B�_g�4 �h.p�0���h��2z��f��ǀ:���n�"p�a��/���7'S0pe��;�Tɷ���i�'�wW��0/�°�W�̡�k�5��EN�b�<�1� P�,��"X�VN�7:�h?���Q2
������f7I�((,)�Q�e�����!��$@�I��F�S�Ƚ��{챪A����&��hUwtu��Ä�L<j)��a��x-��?����G+̟dV�B�.� T�LS�1�Yk��^X���:蠫��
�/�����E$	� L�8h�dXm�����@���ۏe�!�^zi��0BxUz���3�xDe�ri,>�d�0�(��p��������@9�~6t��/�]�2'�9��<��[��E��c�.��D�G��������u�9=��b�&�,���q4MP,�hh��b�I�pp.�3$�)�Ր��6u�Tt���<="�O0yp�{s�8�/���F�`��8��o��fج�t�5�@}>+��XKz�����y�C�pB_Dیmc��ȅQK'�P��|���k&��)����@'O���RK)�����^5���O���7�:�SO=���+b$ZU�D4,��E�����ǈG��X�h��b�a��W�ABha�$��Y�iS��8Q�&�̰����L��,�W�S�\#�c��m���A�,�K�()N֑�f���5"��S�H�A�O8�z�,����D�@s���������/�0�H�H;~)ԀO^��h��Sc���aK�"�!�?L�ɋ>����@�,��P��p��7�FS���s�g"�����G+[����O5K_G� �YYDI'��4�l�w����+�&`5��r�1x�/D����9۪�轹s`e4$E���&Mb�8E�,^VQB��IYs�b�!v.WVqx��C�X͕W^y����e�#xU+nW��T�w-j3���"��������"J�*��Qvb��2��ɇI�@���9Hבu�ڨ��l�2$ȩu{O���~�g�q3��W_*A"m�B|�=2գZ�y��E<q�Y\��`8��By���Ą#���f�/8E�p�t�T�ǂ��Ɂ�8��1s�X�Cz�c��
j��C���=����?�f�"�{����(aL!v4g�:�j>����$:����[^�,�Kx�mǹ|E-H�W�v�m�s�'��[�?�O�`�V�V8�'BD�����!�t�UN�G���4jL_7�u��/4V=�X�Tl�z�ۑ)��u�6���,�H
z��>t�ʲ�p#lC��v��=�	*Lp���H�Zk��#��m�ΩmΫ�a�| @`���g���d�	��a�60�s���� <S䳂BJL��+�9Ɣ���(��Եe�O��w�%�����ӟ�*�9��P�
sQv������$Bi��R��(.�n�d��I�K���#7�ObӖ/0D-&D��wt(�u�F+\f�����^��)kC�֣��QG;&��Hu� v�5S��$΍�zv�0� �h�;���f��BY\�Ftk	�V���L�i� �hUDc ���Pao�N��|k쟫��v�6%���l�F@�X2��'tB�۔iBm���%M�l�2W�P���'�+���>R�Tm+wCQ�T)�v8�8Ʀ`FQ�U��X��歃��a��NA�#h�ii���"ǻ�6�ӫK��׀EUm�[�B�Ƹ�bx�c굚�9p�w�e��75�ү�6w�5F�|�=�(GQ�"�?/CFg���V�%kb���7��U�u]>o`��Z6��)��p;c>��}c��|�����ÚՈ�����˔���tꁚ�<�����vT�5��s;�k>�nS��o����*��U�K�������U�E.�Ui,�K-'�y��7e��.l����(�V'���9Fj����<�\s�5�)��q��{P�;� ���JO:�#��C�/z�j�jk�[��U���N������N��뱱O��$����馛����`�H��)jXm�.�H�T.95&)�'�6�V�%]�խ��X��WSW80<��ε��w��A:�W��wJ�rn��?�_m{WT��\}�՝��O�������L_��5V$���޵Ba��J���κ�I��`O�w�jb��4Q!I���ΏJo��`��c��2%�&����K�2$��"�n�Q"F�'�t,V"VH��(B�ޟ#_uBY���[���ci~^�m�[!a��x'��kX��7(�ɵ#��g�nh�ZD���ٺ9�[����ڽwTM`�M��|n'�Ǥ�?&Qj�L�N>\[{r���ʚ��ʁ�"g��[�u�R��&>� �coƔ�m��|��p�e�г���|G`"z���q��
��R�āzlbS�z���FtBݳ��������&�v��Koy�q��31EP��jы�\��ެ�S��H.�]{r�������.�"�q[L���h�/����B�ݐ�z����Rs���٧�+��ƎjQ���-�6�ҹ�����P���P<} )�+D��
�4�w�Ӵ�,�=?��� k	&��RP>$ {'����a�IS+�����E��n �_]�XJ������� ���_D��cr�I���C\�r;m�甙���s�k��̓_�r�^��3p.X�r}Yq��#��u�C����j�|r�9㹿Y�$Q�������1J9�~�)6�B40��*1��TJ�oB�Z�m8(���9�s��2�2�k"m���!���H�����wE�����:���~c�<�:�9'���<HW�L��l
��q�=sˠW�t��kk�T�#@�՗v2��u�,��5[Tc���Y�c�P�=�-r��q�?�_���j�E�ine�d��)req;~fb.t;x�x�֡Cc��3�k�#"��0�5&w"!*sk=6vVW��y�����(&uN}�S�`�fa�FjF�Eo�) #���|,���)8�|톖~���Tӯ�Ǹ��j��f(������F��r��VH�/�x��&Hy}�����ycG��z�^�v���Ys����?�~�B�eI㏦[)�J���dL��kJ��r��7(S�]/CzLmTb���������u��˼��ƀ,'�Gb��DS�4�1���w���Ѽzz�'��ȣSW��P�3���Qa�3"N멨b&y�PkP�:k�곿5��4��:/z��Uk�[��8[��ԋ4�i�`(�=����n�Őeދ�}���n�_�@�uh��<?�%���i]+.3���@��?)�cg������g���V�w��Iޱ���o\�9b����������1G��3ⁱ�I��˰STs'މ1�x�XJũ�0"�K�)sZd���.&J�j���;$��*BQ����W?.�8� ���>�k-N?2L�����k�`S��u������E���V[�'v5�>�_��׼�T��%�k��B�O�ũ��x[-j��4���2l��N,$�Z���� ���ԗ/4kN�����V�ֹ�1Gu���+T�	�h�h�[�q�"���c�	��04z�&����1�i�e�n�B|Q�枇�b߹����%�߉��'�
�gR�h��F�a�;�}�tf����]�p�9��Ǯ�<�q��X�Nr�����nM(�p`p�Ɩ3��,Tc�8`�v|nR�"�
���[SP,5��{L���5���n�+�p?e,�� f�	oYt�ݣe�=�)8���wE���?׌H�h���V����_;���'���z}���_�s���ƽ��qGb��(��u�_3iRN�W-a�hb�ٯģf��N ���}�	��������9�t�)쯕9� *�������K"lx�w�O���h��΄�'��0��Rc�4QUҿ��[���%�!��m�O�ػ�엦�@��!K?�jf����R�V33ń�;���|��O����W,r �8��'<�adq��������Ž�[M�i�&Zk�%���{&Z��/����I�H��5�K���_�����V��?�:.߄9���V_�W��c�p���턻�jl�t���(�ػ��y��5(�>��w�x�����G�N��]���S�k(k�A]{{m�EnN�*r���_�'S/Џ�'��c���U��8�F��uN2��/��6D#ޡ���h�k��`��I�5�<����BM�i�b��/�՚�� ה����V������ם�Q���U͝�����*�3��4�c���)r��x;����-q+�3�����x^�Q"/\����H�ǝ����z��C��҃Է��g����yٗ�R¢OL�������e�p��F�d�G=��ÚcO���Y��jc+Í�ы�X"Md�����_�h��4���x����d�	�V����֦6K��;�Y��M�j���=�n��p�@�1��M�ZT(�j�����m��0�c��`��ڏ����"D��B��H�=�a��-�@����KRg�n�>R����?f�M>ݻ£"v�;��T�?�J��r���E�*�[fF�i�7_V�*4��9�M}<\� �p�B�PWeN�-r�hg�ǣ�ep7�Y��E��z7Y4ژ!� ?55jٮ�3�s�ū|��?!�R���v�%�ۛ���1"��c�y�UV�>���p;[߷�1 C�����u�[����Ժ���n8�iU�<��D��n勖j���_dhj��|�O<��勖@���x$f�fn�݄��!NN}�E'��N�ڍ�T�,��X���EG�eX>{�|���^��+f��G�/�j�ٻd����N��+�!ye���w�.� O8^!W{���p�e9
�'�B4QO��q~�0�)+"D�R<��I��Ր�M��k4e"qڽ��>uTT�UuYY��8�UM*k�˃���?�H%�܁t�w��5[���"W��k������[��OjK�g�E
E>`���_J����DF�i]3���刢�)�2�R^��s��%F�i�%�����_97�x���k�����yU�6�&G"�o����V.�P�=F��{��0��z������u�� ��2����V�QiD��|-�z0�,��a����B�~�qJ�\�c���(��K�L��Z�rf��֢2����)ˎUٰު�����@:�gu�?�����󌧺����~�nU�a65c��G��ӻ��o��Y�c���ts��zJ�Q���VT�}����;L��ՠF����ˢU"@" �ѐ+�B5��W�������Y+�����[0���{'���=��|}w�̧�3�r	a[�"�zGՕ���x��n�#�:D�h�[6M1S#�M�])���[h��t��V�2��}��	����Z4~�i/�K���vU�\��`�Ա�I�;�iI�u��"��VQ�Z֦ST� 4<�e�:o$�c֡��RL��zE�SB'>���d*/��8�oDo���ټ�O��V.��PS
V�C�����m�u��RpW,���b��(���U�W�ӭ.;ם�T&����e�@�?i����{�2�F�g�ZC�D֨O�Z*1��{z@k*d�x��c�_���Cð�l�����E8`�V��q�4���me�z�Q<[U�Qu"�jW�Z�(�f�������b�vi\�&�:��gN��X�薂"�׮Y��lF���d͐��[Hm%�eo�C�Ԩ+ZF"�ߜ`y�yk�x
.�-iY֚�KFy��-Vb{P��\���g���ׯ�/���g�]��k�UK�>����ty4����o������n
3jA��^�
�=�]4�����̑�k*�f|��2+|���Z=�EwTLb*u�p�J���ݱ�E�3/��s��mM�����N�)���kY�mD��R4?迫=�}��-g\��-���?Z���(b�,5��,�22����6�XʰI}U������C� ��r1lvŌ���ɇc�v���w^�:�w���[�ZfԪn�L�ޛx""B9<t�LjR�	�/�J5����#MR�Y;�C�������猥� ���K��aytr�+�D�5����=���������<Z� V�[�0�h�B�1D���*s�"��o�������ʐ��L3u�;9�ѯs�F����㱎2`2$�p�[��F�ִ�%8Ё����T��i������`.n_�J����,���_���%B&��~�H-f�^�Y�� ���'�}��7�E�Hk%��@��vƩ��ۿ�?!���2r]��@�Uk�1X�2}hn��i�5Y:���ZY�yF,����CY]�d���"�5V����ڹi�»R��3vW���}�4�ASV?|�J�����R5���
)�3����$ VDF ���[��"j0<��0����֖s�5?��zf#T�3�UQ�x������r{E�.�_���J�Ϩ���])����u�ߌq����9昃�(^�A��hF�q l��E�S�՜,=��۲�8U�P�I�_�^*��r�"�����%@�X�[����a�,|&5%��H��Mӫ˰��ȝ%.j���v��F��;��_U�q�*Ɏ��D��0�)��h��SF$��نf�������F)O���Tҥ<ٌ�SF�Z��T��>0 h�^�d45�J�!���eLQ�Җ���+��5��uɃ��ߋ�?sQE)F��a\��i�EƬ�t��y쟪&����s�U��A�c�����^�W*���BL��fV'8�1x�_�P2E��a�x�n`C���H��W��f��T�ժ~v+ C���)[#3�����|K��jh�������dGt[�<�̳�k���ڋW׃�_~����뮻y��u�a�67�}���.��k������;/����}�Y�/�ꫯvB��h.9�7)�b�L�B�+��20a���;３aӹ(��c� ��*�����*t�O������n����x�	f����5�jO����������V[m�u��-����뮻�;�x�]�#�"�����f=��kv�`/��+��⪫�J���=��?��CN:w@��h9 �L�
����J묳��K/�j�ʀZ���{�2(n�߹�o�ZLU��9��L�:��ꄼ��k��	_|�E��8s���	�c�w-��B��^x�{�禛nz��'���`ɭ��f�)��yq�"�,��z���,� F��|ꩧ~��믿��xo��	pX/�=�A�|��+�*�]z��|�Ah���E��@�M�}�^a��|�%��-������k��ӟ�$c��ktl�ߠU34�4i�� ����o���[�y�q��'���·58A4�1`57�`���K
�A�+������8�kz��>)d�Dw�ό>�l��XSx�_B��{>�2ޏ2�t'�w� �,��Gk���ZK-���1Z&D���<,�U��W���aͅ._}��ysQ'�-��, �BE�"l����o�-nU/��2��r�-�,����+tO����-��%��)"��ɓQ5��A�"���@!�v�i�Fuv�����{[Ԃ�de�����^z�%z��曑V�=�~_�̛3<c�W�wm����B�n���-���Oh �w$�'t�8�FC�?�Y�^�/�����Q�=�}�U���1@�o��PF|K�#� �aH����3���>�<���7�x�E]n�7�$�����ӹ�A�5no����SV;�	O���/��T���<��������]��> �DW(4$TB��uF��C"�);T��jF���^�ę��>æs�$+�8���>
C�d'$�%j���m͓BZ�<> >(�~��_�_���E�]}�լ��o�3��<^[��$Bd�̂>�6�c�� �$�&���(I��u1��!�n�*T��D��:�cʊ�ק�~K�(��/�[���q8U?i)*��9�Pd��$�_K��ܹ�z��n7I���`�}���2�ԣ�o�6�	���3�V�M���/�gPpz�����������b%�z���]>�K�7^g���������^����a�~+��a���vگ~�+���SHB�-b�|�]v�s�=YB~	QRV��T:?ꨣ.���gs�@m%���L��X�/~�[o��"�e�^�~��y���.�����T�ୋ9]ar���o#���2�w�yg�}�g^p�H��[�%��B�Ro��v���g�|=庙|�{�1�s��V�y��u���:�[q�o���b�2�R���/J�?���*�.z�v32$��_�_�*�[ ؀�A��s�=��Q�+��7��y���[m����06��nY�m�ݖ�|�߸���aB-D������F�b���/����S�ڡ�������>�l�+eNB({�؄8 �V���?�YY��E�;D�2�,l��-K7t�@���9�a�;��/)��<@��<�4U��!��4�B�����!��m�s9W�>�ՙU��p~].TtM�s���7�d:�����T1�Rw�q]t����q�������~���̩�\`�����������&�|�ng�cM�J���X���/�	VYv��%�^�M���/�
K��x k��6^x�%�ɏ>����?_��|l��Gsբ��[ �#�<#'7��F��8��/��BPc;״I3kNt�o�����>�)\�oρ�����jN9��$K��|o��-J��L>������;�H�
⦼�O�\sͱ�*m囹Jw�dt�������-�؂a�K��mv�}w��y睇Ƀ&�v����'�  ,��Be���o��`E,��~�3)s����nȈc:�e�y�E�`L��=L���;��P�����N��� �����_��t�$7�L	܎za5����V�cHÚ��W�R"��ŷ�P8!�C������{2��?���u��` �G>��H	ޕb�!�s�y�'��*Se��l���<��#�1��ۨ����'p�&�u�O�cY�UW]u��v�c�=�����E���ꪫXY��M==_�;�ybIa����#z@R�S����3΀��;A�rP�)|gO9끕�r�-��g|EEK���x�WN=�T�)�@��a�2a#!�A⫰��)(o�D_&!��������T�Jw0��?_ e��]�8D�7� ɜ~��H���TI�� 8�R�ӟ^{�g˗y�ߘ,���p@�F�p0���7��sk����j���u7�����cƎzG'����/�t�r�]ٞ��G2�_~�/~��x�z��k�jW���߿���o����\"�}�͹M���(���Z�k_��l �㗊�i����9 � O;D4��ݜ���m����CcI�y䩚��A|�{�c�A���"o1�����}�c�g���u���/~�ᇳ��7�p�9c��ԗZ��0�G����jʸ߻c/��W��M7ݔW���ȐY$k���g�%.x����q�"��0T<�)�i�t�.bvD��8`4��	Φ�r�\z8����|�+�PXh`��SJ�t�R������:Wb������}��a����7��ԇ�$��G����E�:)Y)�ќÍ���`^�Z�]�^5! �]�
�n>�����"��T7m,��~���6otKᜌ֎W���
l�(�\%�H�'�tz��8��L�� �rW@-E��i�1ވ�fe1��^ziĲM��yWJ�֊�
�8Ԁc�S�yg9��CK�7�r�"�T�(�_��@��O><-W����A\�S�����K�9��OF���}����7�1C�E,r�a��oƚ6m�v*��Q�G���8c���A#�̄n��1�et.�J9�M{�p;��s�QG/�
�j8l��rS�LAQS�S_)��)Yw�uq�0�_;��)�N��Ѷ*c�8t��u��IP<	����W^Vgq��nH�����S��[l1 8_��Ҙ22^�"��*����w��F�I�֕���Xb	�jJ	i11F�0f\h(��8���.�C�����7�4E��T�u�Y�s�AA�4$6��+��{WnC�}u:��&O����#M��nd�+'�	1�� �i�\1o����S����
�������~�	���sw�B5S�ˋ̞p�	�\r�" ����3������>���^�{�'���@��A�A
8[�j�ն�B�jk���U@��YDf$�$$L	I�<���{��{����~��{+�Z�K��͹���~k��n~��<7:�p�7���"�$�b<�� H^��D��a`ď��Y�X%8��81�p^:`	nW:P-�l�v��q0$����Q�S
o����` ����1^�O�1b	�XNF�c�N=�T���I.�!�5��ڕ�jΐI�����*H(�B���d O�0C�� ,����q����snfW2�_��_a����7wC���'�;��&��R�������SO=ey�������ǬZ�����l�\\�KmJ9�W����4�3�ܾ.s�ڢ�$�v���Yr����*}�S9�ae��ɓ'�}�W�j�{D\i@%QAh�|���6z��G����|E��<lh!���Wf�-����6��4[��C/I�W���0++��Ht1��IҢ晬rgAWH/Ģq�܈��\	*tO�g����=���ᑑF���nVsW)�_N������t�OXpɒ%
`�{�F"�P(���p�Ģ@T՟%�o��ű�{�����gڢ i��\�t��1X��x�,�W\��Q�h���P��}��NsAU��_*g���Rc�fϞ] �!���ὀ�@�ZhWA2�Rce�X�����7������7�'�n�*�ck!9c{������	���ep���J�РJp���֕�w6�\q�Q+|�4-��A�k�����PX�̂O���30���\���)�6����R\,�����M� <���}l�RD�K�v���`ᖙ��Ln�`���!���J���+`E�T��4���x�1`~��L��6�����bi	�H#��%��'ZCϼ�ϛ7Oɓ�G�,"�[p�8�(zL�c]�h%=��c�?������c� �zL���8Fdr� #� n�������N���Tod����w^ux@��گ�z�~?��}�F��)Ӑip�P{��+M?��jy��K���~�e�5�Gqp����ƨ>|]罣�'��oA�3AV=�6o��l�SFk}�[߂y$J��l����s�a���~����3�a3�U��������qp��ywR��LH��U76!K4 �^�������[BX����.��aQ'qK�+���-�~��f2B��LtMg���ﾻ���a$�{�7
?�:q��J�snb 87B�N��4��?�2��� r8a��-�*q��n>�P�lނ����lY����(����Χ<�G�F��0�Ρ+|]���;����a �V��Kp�չXm)����y��ǣ�v4����ICڹ&�ł0gΟy+��+t�Ǵ��"w�MA`^qe��:<�(9Ϯ��x�p����g?+f�$?{C稗K/���)-ښsA��V�)v�a8X=�L�y]��k��M�;;3$*�������|��;b�j���b�ޖR����V�${�����Ԅ	�vZM`�P�����p�%A��C��@8|��l��`��J���?�̇N8a�ܹ�т]�~~qQ�:	jҙ�WK}�Z�����/���_��8�Z����#+�����mj�y������fz��'E�p��@�>zb/'��'-�D�B�9 ��ۿ�[�����+�C?��/}�K��N��K�]l��"�7��(�H��5T�t>���B��-���uk~_"����衇�s�� 2#p?sD���#c'�w'm�}�=��������h��Mm�*H���)��bLbiEΟ�0�1$��_�:�>gΜ�?��=+�Yݎ4M�6����i�,��SA?�~8`���u8e^������5=X�Y>�6�q*X�+���5i���][�]�a���
�'l���OhC�Z� 	i��J� ��E�)������U��A-�5s�!�|��_�ci���\P�T֝u\�b��C�<0�?�AXE����D�~l�[�H@�<�ۄ����ȑC2�C=4�Y򁭂�%2Iɠr��կB�?�Z'�������{�#C�%��+�5����w�_��_2s>���G��" aQ=a;��QG�aAQU%�LN��O�(I8�y&�W���"��!G����UW]��.P\��9����3)s�d)D%1��m����_x�m�46�a�c���k�L�x���*s��c�ҧ>����e3���	���?�#ܮ����\h <
�ˠ�ߚ��g����~6d�ğv^�]P�{�x��n�!�ޠ��� �<P�3y�L�-+�n�X�XL� �'�g1��q�g!�\��h4=�"������zF)"�[g�y�̙3M��"JE[)-%�X�hb�f�;<h�+<Lt��\i���	'���> ��W_���M	^.�]cS�E�^�[�ŦO��u��J�9����R���I�� ��^d��+!�����v����y�W�d��:��A�ӋVV�݂!�
rrRߴuV�v�]�����0-Z��y�9#��1r�ȳ�:�$����1Q2��[�I�*OY�����6/�6$[�yZ�z��,�`��kY�vC�Q�l|m]����C�d�M"��]	dW�KYԿ���tqz���|���f/��$����B:��1~�{ރ��S40�|�� �ڬ���-��a��|�#�ݭ����f�p��-�] �?�+��a+EV�c�Ŵ�&U�����w�}qܟ}��d`�_ORˑG)0�����+MS*@	<%y��ǐ5<��FV�)$�$�\BF�D�$TusTP��(0�Wľ�p�j��H2?c���g�	�l��e��>�h ��{i`ʖ>�Ce��Gq?��s��t��s�����[b�\�ؿ_�b"_� |	�т,�`�X��\� �qx��F�����c�G��5F�U���� ����R����f
+t��-��`�8d [�p�<��n���p�j�+p��+BApV�䓣�d�FNS?��{���k�d	5@R n�h����B��CE������~B�q��a�	�^��fd�f�ߢ8~��N;-�'�R�L|�H���ŝzꩌ�P���pAmEx/H?Xi,a�
BP3r�7`0�}���B�h�}�C ��=��E���jD�^W���r�}��|��ZSEjS�_꼁���.�P�pq�D<3a���'��5w��Xj���>��vY�8$���Z���zY���{�/����-�'����7co��_gAtT����/��t6*�54fYf�@H���FW����{g͚U	�v�{��Xx�(��uJ��%_���A���.%����:Q����w�������F�N���[\t\�����-�j�5��jcA�/�h	�ڨk�SP�O]��.Ψ4KV���]w���NO�>+�k�ب�~E�����)�'$��s�����6��[��V0����m��7�츩�w�GQ�幍9m[��bG/�A��'3�O��'�x"����s~���/�J���$��.��
�z6�m�������������_���p��Q�ΧN�����L�9����ؠ	��Fr���۵��І�� <��0r��e��z 3���,�^˒Y�-	�N������,�ښ�������42C����r�*���1c�hC�X�"��v�I']|��x�n�=����q���c�VE5}����pN�Æ�+ Kb@y<âz�/���9⍪u����;}n0W�+��袋^x���v��Pbv���W��|�Ư�	�t��w���]U_Q.��h�mP��۞{�	1�#&'���-Ԗ��4	���YYY&)2�(~�-�$���)��g��(�Q�ɠ������w��]W^y%4��1zИ Qt���M��Y{�^x��>�	W��4�]w�Pn_�����Ɛ���+V� J�AވG6����Z�K�F�,`H���.� �(��[�����\p��������:A�6W�#���M ��?��K/��T(}����ؖ@h�ł�5_I�y��p ����/���U4$ƀ b�v�y08k��gQ0<�Fh�_#��ů������q��`e+��b�X���=�sT�ͤ5\e������>��66�7n~ײe�,�܂y���' ���0
?��J�1{d�����N;��8��*�@o(��A�͞=[dL�P�u� A�.�������	h����-�c�cƯtO&���`k��g䈒k�t6Gf�q���!��+��0�m���?l F=�	a��b�����!��2$7��[`���$�ڟ���D",�����Ν[�O #+�S
F�f���&/��}���Yٺ.���������GT@�W�1��-ZTw��aE�qW����b;�Ԑ��w�nװ��S��X��v[�4��wܱ`���k���y܎�S��f�EATW�cn��Gy�N����:�!�w��Q�ð/�N�8rDX.�P��`mc���|~�����_��zƵ|P���o-U�d�P�(ڃfn]��^���J����J׿<:�m�2�/�T#_�?�/7��Oe�e�ux�%��8��.���5E
Y����)�L}��I��6V��-�BC�~!`���Q$��vަ[���/�j��O���3'آe�k��@Q���wC���)�3B��@�5${�MZb��P"ipc�~k�K�&y� ���6��K.�dݺu�W'�.q�;Ģ���2�%���lM?��r�w��e���>XMm�ն���	�g�Lf�TP����i^@�.d� /��G����]����(k!�B|��m#�?Ibe�M�V���K�O*�V�ɬ�"sֹ�Z1'lO�C�|n�$Qiaؾ�o��ܚ^�D@p�N�I3D��&�r�u��< n��U_;��V@�$�uF�|ժU�߁	՗�Np�������Ic̬&���`e�@1 S/[�4Blό3�=l�8�e�o��K�^'Kc+@-����W_]w �Po�T�����%_�Y����~���=����ng�wl ~^�;���h��W]�4��n���`�� tT�6�G���i3��/�O�N��HJ3=�r�g���2����l\gB�3u��"��'MRw����y�]w�mͥAFӤI����/��s1󋘀Ѥ���
]�ZV}1�7�0/��_|��AӀ��ʨ��)��W��v�t@����W��ɘ�U�Z}_�1Z�ǈO�����:��Qh�`P`w(�[(���p�	@�3�ev�h���z�sK�����-��.:hz$S�b{�y�RM���1��R��p;�yqů��	��O��mVؚ�Ǝ����s1:/&��z�?���|*��̀˘YBEm�Lw�p٭U]]��UI��V֩Xr�I�c�� �g���--M���Y�-��/��B�B*G>{�/��k�:�P�>��q��1�:�
���A�pߧ����}yUh�iy�ȇ��)�A;�xX��sΉ�����b-�_���-,r����F���-]���	��)�-o�&��[9������|	A�п�(�Mǳv�ygզ�}} ���ȣNE�9�f����[x���T���=��M�P(
U�����s�k��}��6��F�B�4�C:r��=@:�1Y�g�+�X�,+�VJ�k���qt�=�Y%��:��u���������%�l���h`�?�]Aps#K>��m��<�� Cv5r4� ?�|���5�1F��і��.�pA�$��� `�G1���)��(��=����t��\7�L�_�����(��qA�|���	䄇�Q�Ĩ����k�_A�����6�?D׭[�ٸ����X��77�Ӂ�U�	�  ��IDAT"�:4�����-�(8������v@� j� k�F~��֍��TP�U])�A[���y�ԩ�䣏>Z�[p���+u:hS)��*�]m�h'�1/���!{�x}s<���t�Muʰ��{�/
3����lz�3�x�7��L��F:��-�y󇁡�V�3���W�Z�?̜�Ҋ�fl�A��.-	��7&y�Z4����V�'E:+1��Sy�9r0��B��\'�P᷺��AZQT��2h�aȦ�K6�0y�����_�=�&.��.�&^��;���Ç7�����Y��/2L�ůqt�v���=Y^ݞ'6�̡�V+/o�u�ޝ{�%�\I���c�+�RW߸������(7lQ�d!�8����1�ǹR\*�]sIK�����弴��YQ^m��R�?Q�Uk6�,"���E�%�0�q�F"t]���/jb�ʕu`�:�7�y-8�����<4�P�f��a�,Y���*���&�+�{ *zc^�S4Q��A	�V�<
*�����+�Pa�����-�H��C���rڠtp>�O2�k�g���jP�N��V���	@,��-�8�ʪ0_ߛM���ht�ъ|��1����ݬi$�/>���y[�ti�l��<�Rx;�Y@�Tm-8��rd_΋�53���<�Y�Կ�e�����.v\�[l/m �x�N}jݾ3�P��8H�QJC\x��6PM��5kL;Jv CV��wj�t��v2=�rQcc�@m�_��Y��o#_\�p�aoK�
�h�[���c��ZMհ4��-Q�uM�E�*�F�+=��
+$��"C��/�E�o��3��T��]�&��,��V�\�
Öq�R��`��h���6�:H4&o�3p1�;�Mi0�v۱�k<Mt�4�3ܬ�ʒ2rIw����^��6�u1�޵��[5h%+�}t{�s[ w�!��0TF�9�q����A֬�֖�ns/!>�~��C=)h.�:ba�nK�JN#B�\JK(���&J���M�v��;Z�5OC�T!ZޫD��5s�_,�l��B�8_E*�A"�����`um)������]��G��4k����Q�a��ѩT}	��(nk��Ժ����?ѕ�A���ore_1�j�Xv1@�
п~m{I��y� � ��W�+��uk?����ҮB�8X����A��S���C���'-���b��\��v2 g�Ru�MC�]�A)pobV���UY���M�c���I}����!�P�'�e�rU�E��jڢ<��VD��HL�Ð>�g���(���0P<5�Y�~�_ђE-tUmq���6_1dr������i�:�R�\���pA0�y9�d�ds�mֳx[�
��{����ߊZ��'�	8d�P��j�����c��f�XD�h |���AUy(2����	̀����mu��,|�3X�I1 ��,�V��]2�+T�+k���tt�1V�]A�5_�A��y����w)7K�A�+Q*��ʔ�۸�uԮ��S��&�7T�M���.�p!4N�-op�)�n�ȋ�h��'��p�k�ZD>�o��ġ��M�۩�PNm�B\���V@�#�Db�Yӣ�F��w���N��a���l<i^`��Q�k�pg�_ZҘ���E(Fb^h#��B[�p�V����)�[���xs���&�S_Q@^Ƭ2>͘�5�4��E�R�i���T	�bcdo���d�S|�(�Җ��ֿ`C\x���ֶ��Z��	���r}�����\Q�R��)���=),Vӗ �;�0~ic�ucWO_��F�kIkq
�w�(�l ��o�4!BȗBZ�d]2>`���_]�ͩ���mK��]C��>X!�$��+n�b׬Y�~�zSp�0$o�yc��^�f�WJV�!n8w/��l�2��%� =+�DϫV�*���Ɵ�ܸq��׹ߥ1�իW�JHlh2y5��
�XS���.�⇶Gj4C���j�C�$x���*Ӱ6�	}T�t�[����]b�p��yL�f�6��j6VW�]y網!ç���p����h��v�x<�Z��tn�@�}�u�ts�a��T�
�./v�L����=7ʑ�ދ���3�!LA<��I��4ѻ ��Zonsy2i�g��M?�a�ס6��]�ָ�i^8\G}b�>	*�66��Ֆ���Sӄ% Qh��g4��m6���έt�u}�~�]q�ڀ�m���'4���:#G�l�)a��V��j���?��>k|���
lI.�����pP=f���[ݪ{A��̊ �4@x<����0mX�dK=��"���([���fA�ѓ���-�A/�~ޒWȄ�-�ɫ��Z��=�^oR�b|�����9�B|�R�v��0?��B2u������#\���K,H�������"�l!Zh[[(���
v��%K�i�����vA��lVa� :�ڻ�o����M�:u]P�5�E�f������ d��8=��#�!B��3׽~}~Y}[F~�=���&�Z�~���*�}�G�c��4n����S5�D���C����Gh����O�q���߾Y��?�l���@jP�&۳:o��o��[V%��
5��V9GW>\����HK��͛7�������E��H�6נ��x��f��-mIԶ�AL�Ϊ9��J�<0q��b�^�%M�v9U!�,��%����@��ͮa7�Y3���m�X��50fV5�S�uM���o~cw�ؽ!V��߲��ʤ��M4"k�^��-]�ԬE�t�%�#�lAF����o9��L���<��ѣGې�5
JUap�I��A����'A��f7p%ePue�Bo0�H��,Xp�I'A=A(3��H�P.�34��+*����y��;e�^ǅ���+�'��~���;>�¨^�O�o�&|bI��K�:A�a�0�*v�3�"�<��S�,���s8.WY�_ŗB%���ЀR��<Y�U}�BG~��.��w�ä7�1�a����ɓ'7�sc�p
��'S�33q��a��ٳgG>5�x���%��-��{�F�B�6�͢�b�]DF�h�o�	�l��v��6��D�B0��4lz�K�-�� �K_|�E�^�ћ���bY{�7]:����;ҊQ.��������vՃ��fS�L�h��u�#R�v�I�[g��Ǣ����s��$�(: �2'���z� �[#Q�.ܝs�.�jF�17�X�>�=f��ּ��B���^�5ZÜDɖ�#��U�8<�^�W�?��r��>o���+^y�����8��}.\�<��=Y^��PdDKW��z6k�z�*i��K�P���Jݛ6�ow��dHGwT*w��j��^���l��KK�+Eq�����_y橧�>�X�����W�����t�w�u�-ai���'���u��:4��<�F|��G!���\�wD'�=�؉'���k���e��k����?�����1?��~���$�W�-g��Pw�}w�#7�`�Óhy��Pi�.P����Zpd�̝;ׂ7�٩���{�v�i��y�_\o�-Q�n�
 �ka����Y���֏?���{�Y����4Ɲ���㌕z+Q��}]]w�qg�R5��Q��d�e���Z���?���GqTK����j��u5�\R�F�lJ�<G
�2���nd6�б��]+^�+�$8A�(�\Dl	 }�m���8�j�ޖ����{�ע)��o��|x�GxL��3O�dt�4[\h�h���:��'��*)?�j����K���� y�V�?��s���y督�ԦLm�>�v�n��v�z��#1DF��3f�(��6f��\G:g�B��m���"�E��S��)�ܬo��o��J�=:[t`ĬY������+�u���T83��	�1���v�<
-���b<���C
��;�a۝�Jذ�׿y��Ə��z1�1��m�I���;˗���s�&O���@������q���?ё��s�=��S*�m����N@��~=	�*��BX�rه!�}�������x�裏5j��aP�[��>d�(�a���HH�����ci���8����������oJ��hL����CG"��x��m�9#��#����U��ziJG�/�S N�"��j�P<�w��Ο�Ҙ��g�*���w�y��u1z* ī��G���q�����n7:o_B��'�����WǊ~n�����sW�{�D
��G[�v}ې��LR�:�	g'j}��4i�P=	`eO8�I�&�>4�^�f��) j�2�/�+�؞{�wY���à�� +��_�JY��+C#��o��v�i'���ц�)U{��Q	:�rl�Q�h!U@6]Z�u �+�ӹ��`6��Q@����t�d���a����q�5ۖ��M���[n�����fEX�:*��Qf���_*�!���6X�	Ao�օ9���(����}YK���-����l��Nǒ@������h��~^�nG}���Y�tKkH_S��k�#\���2O��P�j�T�֬�ɡ%�*p%,��,ߣP��5i�	b>��O�*\��ø�!%�%�5W��ӀJ�_=���0.��^!�	p��b�/���}��j�8��w9a�t)��z� c&���7߬�r#�>݊�Or�����\/,�HА/a;]S�7!��c�<ðQ��i\�Q���y*B���j����]�|���a��n�3����
D"���W��-��#����7��=I��cea�\��޶ֶ�l��[�:�;�,e8m��q����fc_{A>�i�U>��J��[͢�k2�t�>����x��*V�R	�f�'~��_�����֨T?�g =�m;����#I��RP&rڌ8�#�ʍ7�x衇�7�.�6w.�{�R����;K��k�=��ȗ-[v�7|�T�������B�7nT):�=u/z�� 0��C	Ip�A�C�S��8�C-8�F�������c�=v��ԨCY8��8_Dj�&�db�|�9�%��=_*��٫%_TW9����.��Ѻ�Xp���w�q�6eL6uw!5I����]�2.;��K3��!~����kF|�x�bx��N�Y�:�g��Q=� ����ȱ���g�JY�
]q6
N�J1_�oT��<mC�'�SN9�Dy�>�ל��MmV��·ز�s�����l"O�뮻��ӧ��`���,�2�M7�T�{ɋ�Dw�}76Qe�,L��4R���ISq:0�f#�O��=�y�n4��,���L�޾t��+��B�_��~����>(&x�S�_�`�v2LXmtl��%�c�D�혵�[Y� j<]]�Pb�b٬���}�h��2�Z�-n`�θ(ɳC����n�-���A��>���g����1�I������˖�l��R��_�jP��s�[4��ET��s��di� �o=��M���ꫯ>묳����*�۲��_\6�3hH��0��5i8Çr�qc�f�>�M�P�gȊ���a�PA����������^�2A����E��6-
���5I��=��e�u�B�{f����3��E=���2��L줻���Z�ퟎ�ұ⍝��Ī��v�ԓĵ�I�r�����x*�n��|�4Wp�;?�[�1 �믵'��W^y�U��G)8��,��{����;� ��d���RV������ި��Ud$pϏ~����5���.x���~jho���'�g�q�GZ�3��� �fM}��\ �[�"_��@�`h�*s8<(��|\;y衇~�ӟ�Y�&��4E�P�O�_~9��l6�{��Y���+Ui[�?Q=@���-9't����^{�g>��m�io.��RT����6ĥ�+/:����t����=���8�]5Rn����
���/N<�ؽ߲?�)�Oj��!�rf(�\v.��5�u�f^M�Z�}���A.�H�}�:>1*iYQ=��?�mo{[��딞!!������[�/�"�ꪫ��g ��!nׂ�6�h�d�~``B����$�<Ez�8��3�-� I�|r�?{ N.<���X#�3<�<����E��h��!<m����pZck�4Bd{��n�!��lZ�|^����0*J��hbc)k˗/��@Di(bg�]���`[���nO��r]�\S}���rZt��κ�?q�HA��u��j��萗�ƿ�]��5��B(�����dE�ϯ�r��׵7�z�V?ξ���݀�V{����c�;�NT�#8������/ߥtU�-Te��Q�%6�n��O~�b�z��H&w��f��v�Te����nge�K���%�(fy���\#x20;N���H����lv����0�&�\r	+����-�)8��Ah�O<q���Sa��e1�[���PVޠ�A�5�:U��5�F^T���ƅ ɮdr��:GK`?�яF��j��4Y��y[�U��_|�Ÿ[�{z�@:|�SO=����i��Ec¨�l��^4<��.�oʳ Ġ�3}�z��>��Ø�3���F�?�%t�2����V�^[�
��.��Es��S�Ni-�@�����p-P�
d����0�=hC��?��s�9+@�J5`�d�Zv����Oˡ5=�|)��c��#�8B(����\�GDk-"����i�j�!4�*f����J�����'@����� (I��2�0t���^z�.�������l�-��ؘS����*)�ͅ���cж@�6�����~�3��x�\|�!����� ��p�E���������s�U��p$���f���ltY��e�����ᶶ�.g�  ��ʥr�֯)����N�hE���:�}
��8��LQ�Xi���������MNl�FaK�%�q*��4J��X�0�{�����y�2n(P �#��{��UHf>4�Z~�w��ɓ'c~��:O�Ӑ��OXfh\��k�!U�={6À,v��9�vn���1�s�PO�`R��i��6Љ�E�+GI��ж�^�c�.�ۘ�f?�袋�$aK
U~-��g<V���.���^��G����q������?������ӧ�*�R殾�����iWM�ƴ������Ժ���ʋ��?�=��;��_�j��F�vV
�I&;����������@ �6�lcƬ��c�"���T�h�+%:G���?��v�qG<R�?3���-[�'h��`��İ�[��9�쳑����C͟��H�*���+���S��0����7��Mh����#_5EB�waV�Gy���l}�Ǡ�<�@zf��+u��ܣ�>
�K.��n�p��I����� ��.���1=V��W����!}�c[rNb�b�|�v�ܹ������ĉ�|��̕�}��%��˖-�c���tI�@<h���|��YY0��I�2i�#,U��(��K!)�%�2�9�r�=T���G��e��|x��&�`I��\���W\��N;��Z+�-0!������;�d0�l���}C��id�$+����ɑ��@���a�4�2}�ס�e˞y��+k�5��4�b��
j���/ù�M�ɓx���O~�bݚ/W"cd���!�������un��ַ����������J�Q/�p�-�7��P�\����̘1�eYsR,ad�����_��P#c�����/���M��VP��p�S �jА�_}�0�H,��O2�/|�L ��c��ᝇ�h!���p��r��j0z�8���&�P��F:'
Rb����/���|#�hhʇE"��կ�gpGky����1w��p�n�֥�Ѿ_�p�d���u
����h��<�s櫯�J��i]X��#|�ˊ����W�:�b�ql��ͯ������OШ�뽨S���O�z)ȥǴ��Qf���)^G-�����y�{-hxlI��k�04�ci�
��ӑI���v�kS��'qex+��'7I-]����:;�[�Z�Ҿ���B��˒�3X����ʗ�E����|�_�q�W���2O�U���tr1񍉡�����FkB�M�`�� `T�������޹<�'Q��99���E��ظV(,��*�0�z����?�y�ϬT3�MJ����|��N�2Eq&3l2���9��L��NB��Ռ� <4���?�:B1KC~z��"����S���] ����p���_��׾5�ï�j3B�*,��>(˚緤�Ÿ�+�CL��ۿ�2	U��r!���j��JvM2f��[n��w��z�jӡ�e�Բ-1į��ʼ�%j��T��o��<a�{�v�c
�4gC�8u��J��pL>�]���s���k	 Y�3��k��$I��c�|~r�m�!�8 �'A�w�Q�R�U���Wِ$�zl�XDy �,ķ�yK>���6���΂s̅�W�	�q�n���_��_ �I'�� se�m`
�%+�.^��8Zf����gA-�-����-��սlP���o|������$�<��ː��[�֘M�K�\�/~��rK��z�1�������~��]l��-��y���?��EՏ�é8������7�r��K���G�;���*� ���K�m���BZ!#�N�5r� K�25$���9�lF2 -��;[bt���ԕ�S=��Sp+ˋ��\h�K����z).�two����"�u�(�bp�vt;��I�����#1�	 ��S��oY���� '�ls�ǆ#zR�Q�O�p�:t^�U8l�`�
�X �i����Z�NV�A!�k����D��F8f�jP1h`ET�u�9�uh�dk�M�B��B1#������/�bf^^�=�'�kA�5�����5j�A��*�S�Z�R��d�8BLPW2+�a�a֭����):��K-�oa�1��1h3�͚5P���IP�KZZҍB�-0�qi-	T�@:ɟ�I�<9���l3.�y���
^��v�W
����u!��(���/A�vub~�2���h�9s�@|�W���4�C�O��L��aq�.L0-�'�@w��`�5k֘?c��n j%�#CT%�U��B-�_"8}�'�����������ˏ���01I!i�'(�����/�T���?<�c��ĺ�] ��z�ҥ���Y�Q�@������v�I�J�c�J�yӞ�R��^��!�u�l�+7d?��^Ko&޵��#��k˯�1Ìc�n�ՏNFk�b�ʑ/�,��W-=h�4���<�:ǂ"����m<��q���{����f�P�V삣�``�Ї�v�H��x�M7����mh� Zl�������?=��x)0� 9��������jP��D�4Hm�u�5��M��c��[o���K/�������E7�c_�����eN9�3f�O26�=�#,�u�]w�y灇\nť����hh�����?��O��_�FH#�m)�t�d#;C�kW�����n6Z�,�E�jնֶ޾^��٥�>�O��^�G��Tk��T�L�zk�!��y�!4ȍ7ߜ���f�Z}s�dDa6��}�{�B�	O���H��?�9��cr��"윮����O�Ua�<0N��%��G}����`j�S&��(�/�i�����9j�=�y����ֳ6���0�y��IA����c�n��'>�O}
m8b�sm`Ёy���<ZǍ�6���/F��ӟ֙�R����/jx(_Y��ՃrM�{Z�#��a;�<�HPK(z�Z�\�O%K��v1����������˻���:���U�������袋 O��3�Omo����pL��~�덊�
��1lz��k	f�W5#>�>Ͳ������_��_u��y�l1�����ٳg_yU����p�t̳���o~󛨚�~����3�4S�C�A|��p�����$�BoqpJ���J����9�2�og��󱙻b��K�-5�gH WV=6r��0%w�g�=C��ׂ��>���r���3CB��;��q�\�U�Ё���o��v%��~[�nPF_��zfQR$N�72�*�5��e���7�Rҹ��LW8�F��&ջt/�3T`o�N젔��x衇�;V)a��QI��' �&�5�w��'~7^bu��7�jPeGqİa��ʂ0 ��e<\p�T�k���1T��x�g>���9����#�(�q,�Y�!h�rW�@+ ~8��3��'�p�.��T��/{� 4���9�ۅ��&[:�H�������~��'��Qp
%��a؋���
Ɠ�;�����*� �兘.��r�$l�n	��jKG�A���y����^,&R���<��s�3 �}��G�Qɖ�w��Bj��ܹs�
п�Y����0q�D;�&��Ap<�s�9���X�݀�fw ���g>󙷾���ӱ����_7t˵�^�aM���AC 喴��u�T#WuCz�T���g�������B�绺Qղ����ҚK�3�E|�O���Ҥ��DY`�N=��C9��^���Ƽ	Jւ)6+�
��;X-z`	�߰�������@V��P�?��OU2�x� �oIؐ����vw����u�]M��t��!�fK�/Z�f���P����O1'�x"HnҤI���Čp�,X`��BH�Pw>�Z�����g?�4�B��~�ᰈ�7��B�
uk�ׂ���b3��reB}&~R���cۆc�`,:�2I��^w/[��	�Тz�f�B"��;���N�*�瞝s��w���s�d&ٞ�ˏ��\�����_3^��0�|߇���^�$7�x��/�e):�����G��������S��v���^�X��\����z���u���eE�C|�e\�$H,d��.�y�雐J.%�>��i�}����/�.a�&���F|E]�n�J��!����X���{����@��;i��-̃�����Ђ�-��cQ��H�QG������p���p#�?��#�|C� �o!%�AN� 04��.>��q�!8"�Bx���J\�Qqad�k_� WK���u�E�k��	���%��j��m������1c�(���%1$��E�G{��'A▽���������ϰ�b�� ���&/�����RεJ6qWk���s}�9/s��07vmڴ��{�y�'N8�$f�?~�xu͚u,:��>��li	��ݚ�|n���b �

3��̙31�����_��-'��pQ],Clc�" 2:��vu6T�pYq�m�s8���N�!u�Ca������m�#�C(j�� �)<�V�˸.�t�P�J�i�^ ,��S��w�k���W ��@��x���<�m�kgI!�Z~��C t�r��w4�4 ���AZ�Pꓑ�r��O+3L�N`i���"@ ��YP�����ӗ_e �h�(�P/�Ɣ�-|�I����������e,�xPޚ��y ���o��Q��`�xM�sP�gf�ؙEjk�buW����g�J��/����=��Ϝt�ɨ�P��v�9���4������)uo���F��w��8 ʒ��k�#J)KP��JG�'��\��G�I����E�Q&騡V�xp{%�MU�[vIÐ���w��b5�t�۲��-w䍕���i(�6�PN�����7�*{�1u>�� b)�	��&I�9�؉1k_���~���
����K!�e?ڔ�-b$��?+�u8�3����;��<�@�虵��h��OK6��+�#�ΡB N�,L%�VM2�[j�3X�0���е���#���V��$]�lb�g	�7n� >����6�$&��H0�h{O<�RV~3�/\���/f���2<�B�!튋�H}�I5�ǟx��ێΕP�2Z�d	#���_&0T�EH�u����
��,�`��j�U�j���}$�n`�M�qg�O$z�n6JD*x�ʕh����c�%1�Ѳ�"WB���0ۉ�mY�P�[��b�a*K8�VI���] �4���'�n�ԍ�6��yc�[n�Ӵ�|	�<���ȫ�J).U�4���j�Iw'm��3f��6��?��y�����f�:�y��Y�xы�ʥ<���?т���4R���|1>A�իW�s"�@�μi��ee"������rƉ�-�!H�<Ht+�WpN*��q'�ܜ�$H	�5U]P���<l)v��-@Մ	�5�D ����mx�@UY�2��+�h�	�������x5���)�(+���8���^x!������9�������E�
v��)�4��ڨ� ����9��ԳFR�g����,h��Oh�������?��'����*����ۆ�mX҂m,Ȫɢ3 ���.��Z�K�$�4'�i�H"/Z�f~�͖�\�5Y x�tC��m`d�Y�j�2aZ�Ca�?
	R��l	�ʽ䷌�G?���Ӕ�)�Hdi�1��E�~���|��Y�f1H�=��2�����󨤁�u�O�}�Af��O$36y��P:W���̡q*�j�\3�W��
�p�Ո?�MtaÀ�Pe�w��*�w�)�,��Yg�5m�4DI��������,��l����#Q��d�:3ƗH(3��-Ä)Q�I�?l�:,()V�ɫ��c�z��V�z�����>�V���K� �8��,P��%�+�1,����?��-Ojp�S"Ý����{�t�%R��^{�u��uЇ��v0�<T+^�ؗEQ�����3l:M��_˿�S'�N���(�ː^b�ÍS��6:5'tg�vY�	�i�iL��c�Y+��sh՗���ˉ2�d�!� 4~�B���o�[�йnfE�T.Lt��L��@��x��E?��0I@zf�h :��-�� @�u�GJ��/Z����$�ɁՔ�_�Oe澮�K�Zy�k˶�*}�k:]�{kOv�o�g֢�|��zKQ�VI�̢�F���������ޒ��1�OB,�[�|+��Q:sې�_ø�6������)c�0����|({��س&�*o�
����p.uxZ?��P��f����{��R�����������p+ �����X�nu���9�,��"�D�96/�Z+�J���û�2�����6��G�7c��2��21hIk��]���e�.]�6�����ܧK]]i�ԇ�)�]-s$����~ �u,i�Sa�OƓi~Qq�ʚ��g�󠬨��֬��8_]|�.o$�9z.o���5���F�q[��F�A�gazYe�K���+���y϶x��ۻ�I3`E��K�p�&��4�Fkrtp�)"S�6��xX?r̈́(+�P���f�����y\\����nW,�<LcVB7���0�����d�pl!o�1�W���l�j�] }������5G�ڳ-�4ޠ~_�	�"o���1I��P��F=��;o�S׌Ÿ�7d�j^P���|xB�m�ޅ�j�����p�z��N�y���vn�Y��P�8�Q��A%8����D�<�[��̡3>����N��gg1�R)�g��V6��[4���M�5oK���_����p����#u�=R���I�v�6$`�y�a
�V<\z�a��{�"�y���g�%X��{W��T�}�f��D��n��:��K��f�����������.�@�[��yȵ[4<���4(:X'��Inm[[����tqD����%�Zz%ɭ�p}�z�qЁ�8��׶D8?��CƎ;��Ǳ��k��9s�3���=�\k[[~9X-��/J�pe��۟�������2���\v0&�O��h]_��hʔ){�e�!#G�7j(��qL������4�s����jk���GQê���qdnF�С���̙3�kR�!Mcǎ�={��9sZZJ����V\5��OH��?M��C�!Y�ûJ#{Z��q�Wco�f���W�/��QVn��Tˮ8������M�R�n5[���nl����a�jv�n�e�⚺��v����Qo;��.)�^������*�����Y�������5f����Q3��~q~_9rլ`PK���[J%���w�����O��Z�9��I���k��" �Q�F����Ƥғ�P�蜶����7�H��A���"�Qp�I�Wnk���O�7NZ�������fytY�4��0����ӧOW�8ɚ<y���g�_ink������Z5ml��.(������ۣT�í�ҭ��iM��S1X��(?���25�V>����cȸ1�֭�r��cǎՆ@����m���DK����/��۸v�������(���6~����]^���x������k���ɟ�(d6i����f"�t���yr�m��Q�]v�e��ź��6�X��ڶ�?ۖ�g{��A��]��!Y	���,�^eu*���}Ĉ<9z�������FvZ[K�}�V���Z�7m�sC�.�m�k�UMֶf7�TK�Ua���K-�//�4z��4J[��Tri���h�� �-����LZ�����������Y���	f�QQ\����,G�\j�s��M�1c�c��f�m*#;W�^=����.}|�O<�0%+�=s�СC�:���y��s��Y����+WT�������0e݊�\^�V͊���Z)�����7���4��1qxSZ���:�zz+����g���n��umm�I��Çoܸq�s��)ǥg�9꘣u�t�ĉ6lȎ��h緹lr�R~k�#��)y��H���7m�6dҤI;��؉�t�</�����+g͚�ڒ%��]w�u����'� �{{k�ev[����l���n��,��ܙ�n��4�J�ť$?�X�˰�`�������(no"[�A���7�7����GVRI��s�"Q�T�f�T(�>������{7-]�bţ�>����\���Q�^{��ٴi��f��⋮/]�d��m'����;v�СnmWN�?�\ެ���O��?�,�ZӰ��?�e�\תY��裏VA���DM� 8�-���բ�4>���U�ӦM{�W�2Gq��xy���C-8~�����X9�c�?����-&I��w�a��w�yذa]=�*GN�]� ,_���E��ϟ?}���%��h���Ņ]]�i��o���>��%r궀D�����zg��&�mr���\��ѱiTv�=�Ӽ�o^���E?d�伨^-�JyD?�Ҽ"g^��mQ~>3�4��S"����f��f�-���^�!
�Zo��[���J�����YM�,G��:l�v;�=۶��1z��+@��*}��E_ye��J��^ֹM��Vv�5a膞�}����W_r=i��e�	+&L��:���8}ճ�]O����n�c�[�c��Y�7���>�d����K_<�7W'4{�w�����3ob�$�մ�3B=|Ըm��v��f�aKe�uȳ��#F����U��ZZ��z{���ܼ��1|��1�L�
|)�п��k��`���wko���?������=9�����п��;�?C�]]S&O�n��\�>���Q���OuSl���U�ΡÓZe�ڵ�^X��t��ɯ��RVR.ތ��=������Ǜ�o���Cۻ7e���m�O�O=���ի�tfUS�Q��r�{Bu̘Qk�6�~��G��[xt7A�_����%���=Z�n��sw��h-��ip]Λ��I��_jmM����i�v�m�R�:nܸt��e˖���ߌ�c�m��E�s��７�Z�ܹsۧ��ݷ��]��l�ĉ_X���q#��5��N���W�y��߬	��|����?g���&���O,�{�'L��Ғ]h?|��ٴgf]~�OA�k֬QŒ1cƨ*���Z�ڑ8�?�4s��ŋoڰ��k�S��~�O
?�[�������_��s��o���$8����k^G|��o��c�&��?;:;7m��N�y�Ρ�ٟ�E�]I:8F�R�������&�諼Y�s����#�C�{�WWmqCF����ޕ��Q)�����KƏ�1}x�Z������)��jQ��Z㴥�K���+;.��V��@�۬"K���3�׽J�=��-���5��1�<��G���~�Ŕ�U��[�
(��䠇?׵�})�U~#%M�_{a��_E��q�2��B���>�^��O7�q�S��p��q�,��z2]��t������)ŬGv)����'����w���:�x&��qvI���ik��R�d7Dd���?��v�c%뺽��io�v���GTbW���{$�4�,�[JɄ�C�L阾,Tٶvڴ�t��M�F����W�r��W�.X?n������c��Oo۸���[׭OW��^�1���-un���W_s�n/]+�]��e؈Z���֥�]%��Y�j\R�O����\���墤Q/\��f���-�nJÈ��1�����l���e"����i^�7���ծi���٥�&D��Y�)��!O�Bp���1v���H��Z�l޺��f�W(ב�!R�Uyb������]�ͩ��H��6��]�j$�M@v%�h�3�d��mE++nbnO�_x��VEl���LA�U�3��Ŏ�J�Qv@%�
�d�@�t)�(]��(TY<ͪf�I!��Z��K�L�0�Z��{{W���=���Z��1��s�W+o;i��/-Bd�����W_^��̝{��F�6y����}���tq�)@a�{"SW�k�4xc����&j���_ʋ��T�]R�%06��!����Ç���]�Bu��]�*U-����ܱ���#�:.�;hm�F�~B3TLg�72��ɮ�Ӓ9_a]Ba�פ\a3�o�(���ZB�jT5&\�צ]]?���\f-R��d��ͮ�O�>gG��4˥r-/u�_��XI6�L}�*��pKN�jM���W��\ە��4�=�Λ�f��_�z�ǎ_s��cF5����+���Z�~ɊU3G�d4{���{�'��d̓���L󈀩��k��P�k�lA����F�P�턆LL��N�&�î�qѠ�4V׺�^Ջ�I��.��S��Z�:fi�悻����պ��$��f/�w=�O���_��њ��6%\�f����E�u�5�B.�{|�[�] �2jL�>���j]�	�6�aÆm��Fi�����=ٕ�؄F�IF�a*&�������Tj�j}��r��oܯƠw�qG_匮[�.�"���5��7��;tEV1h^�}ĤI���f͚�_]w@�ģ��(�d�L���6�t�d~o_��826��Woܸ�Y�v_�iC3~5q��q�����kתs�����u~E��Oa�*�O�	��%��ׯ7Mtͧ�+�qX��%�e2����L՚�����cǲ��޾իW���k��P���-���A���_�����TJ6+�j���˰L{[;Þ0q,�.x)�����ΐhu[;X�r%+5~�aLa|��u�u�Q��7l�m��-x~�=�x��GH����m���3g�d!E����\�zZ��|�>��]�z��::z7eNl��dʄ�@���5��L���2��#G��λX���֡3lW&K[i����y�
�Y�!�9=�Pݛ���=��mtǰ�'\h{�x��dY��3f<�3t��M>��:݊Z J��y����}�M�leG��_W�X�(�D=`�u����v�Qn\�M�X����^L����>��,�F�J�kd���x���_S���HUk�ښ��h�$M�#��9��x�b����w��#ξ�y3�i��i�e^fG�с��N������C�����7u�Ut�=����{n�6���n�ͮ�K����x<̒�^٫�>D��K�-}饗2�U�L������ȑ��n���Qc!��%�˜wOLC��u�%t�� o��H�A��ʗAf5��U���n��8��O�?<�z�<y2/��A�_&��9ǳx�n�5C����d:D�3�CF��L�-fޗ���ɷw	�ޱ��>�gt����g��|fןߕ��=	�-�%�K��HH	��l�o! ޢ+�uO0���Ԝ7�'�b�f�:1���)�\h2zt&��Qs���y�!���Z����,í/˼Ϟ�C��+�˹2����a]����w.�twϝ;w�}���f��p�+y��-�V"�,�N;�,�j3�K%��ޠ�ԩS�s�K!O
�,Y���u+6Ԗ�4W� D�?��q�0��1�#��]\�%˹���@gT�*l�*���'����_n�֨�0��MXdY��A|��8>m#{�����U�d�Ev����M���. yR���V�ނ���C����YV�)@xU �,^Ь�P��5p��W�! �a�⊲��6^ W6elF�y�ۤ���Ro���9>C~}Yy��׽�i-��e��-q�����b��y����-�q�7���ׇ�>��N:餽��[�l� �q�7�}�݀ ��K7H��7��e;�Î:ꨝw��!�� `�fͺ��;q���.0*͈���-nͪcގ>��w����ȷ�>�����r�.|v��5�LNc3&���b��8�<��X-���?A��~d^z�y�F�Hǟ<Fo��߻��.��bp�SO=u���?��˗/�âLgG�LJ���^Ϛ��}�q���P��3$������v�m�}ú�2�ot��e@�F�>i�\햓R[k��UG��̝�9昷z0J$>�1�����/�ސ�?yɺu�׍��=�u�;l���kG��n�k��M���=.^�<ӡ-@�am���Z�έ۸a����ː�{���=���D��N�=g��0��O<��|��uk�b��+i�¢��X��HA
�Z��⢤v�}��O>��o}+�
�w��u�u��~����"uפ۵J�c�{z��2�?����v	�$�̳�t>g��DM����!ί|�'g̘�(����Hx�ѭ����s�).�Yܯ���(,�CB�C=4K��wN�4���F�
�(o����>��O<g�@[�Z<��PQ�NT �n}o��.��Kt��r]�!��G�����
�ʌ	Ձ9I�AO�2lΰ�	�.�����{���^2fWY$}��P�_���Q�]�&95 Oe06{��	'������r`Ԗ9-K�>���,(z?`H{��8a�R2�����c*�!��!m}�JG�з���G�k�n���rˢ_9j8�������1T
sh�p޵fMv��;��;^}�e�Aꌨټ�o�)&'�z�{�C2�<���8��7����I�YW���d����J�㎃g%A�C��~��,X �^�j���Ĩ2�2�4h����v�:��1���B�!W�4�4}�~�Yab�oV�a�{�'�ė�H1{��o�nR��sxꚨmr�6�Ř�o䍋-z��gaHȮ�b_��h⠝�\��LczꩧbL�}�Zh��s>���G���FUjU����0�w�����r� PY7�t�=c��߃R1~�o����1o8({�����Z��j��z$:� �H�b�ZV���\C�~�r�.��3W�\��:����2�Y��?zĈ!-�	�a�y-��kVW{{Əݵa�駞�ۮ;gu�ƎUt �١� �4�ز�H��i⯳�LC�$��*��~�C�ca@��Z\�C!C3��F�{��)��B#�9&	ݎ�ҕ���k�F�-��~����-oy��?��@��m���Z�ͻB�޶���P���Qv�G��@w�<��Ō2l:gH�� ԩ	��6��'�H�Gq�";�:`8P/���Sj1�A�4��?�5.��p�)���L�N�����9�XEc��Q��/A�N� U������z�mv4�ڹi�F�G �y����X]�$i�$�L�W�KZ�m�j���O�Ń��a�h�2������v����.��Tjт����?��#*hX�o���5 ��_��_E�o�G漧k��g��~�=�y0H+g��|�ן����^z):]�8�p�s]�.�"�V;��3e�ֵ���}��vĻ�袋��`S�P�1�h���;��ο����>dDM�v�el����C!ZWrX�[�a��S�On>�>����˿�~�X �g}��ȣ�����]}�՗^�y��9oh��7K`�`{ݕ�Z�V��8y��}�s�s<�kٸ���%[�%q� �������w��^[>���'����r�_>eֲE�ܒ%��.�X�hY2I�Ŀ�jOK�����ţ�������a�)��u��ÿy�.����2Z��J�O��7�*ܿ��9s]r��pCBP(�_���_~���!�:h�?Ŵ���ʺ�j�I���YE�\y�=�Pk�hG8�.�1P���uN��ZX���G?��_��W����)`���&Ӣ�>8��"#SگSL��яx2���'�=��_��7��ػP�C�!B�;q�t��'�K{�o�ۏ?�xv�	��s	�u�����>����)� ��;� �  D�òM"�Un�ZWdgA!�'?�Il�ն�V�ϐ#�E%~�{����pC��b�h��,�Y����/��<�z�9s���_���6�s�=��s�v��w���>�+u���k7NӞ�7��99Ӳ�Y0B
ӣ����	�i��X�C;<��kⲓ6���C��G>r�E����>��M�� 	�~����g�OV�7Ё<��<�Ә��矏6 5���oӴ�����>��X0��$���)9�C�k���K.ɪ�5DF��L1~���s���
��g=�t�+��nX\q�?��O���}��q),bǻ�p�Y&�Oq����SO�s�9�D6� ��#Ptr�g�� rj!0B����`����8E2���P|��!Gȩ�H�������,oګwA�U������s�[#�؅?���Dp1C�@UGy5ի�C���,�TG��H4�Ў�b�$;�;|�T����ջ��ᙎ)���u9�gpb�O�fX�t)~��h������$r4lh���|��:n���۱�,�����(������
!�!V��p���c�#�������ƄR��@�%�E�Wav�!J�B� 3� -Ɯ|�k�OfQ������B�DR�x�cL�~��ᨇ�S<�ҙᖣ�\�+8�0<��,�)pi ��_��n�Nq�:�&�b:_��tȫ����v�h �#ܮ�s�D�9�x��gc#���OJ���O>��Vd����<LVxۺfQns-���R�ť��Z�%�-U� ��R���I�D����7�������.o�t�}!	!$$D@E�A�A�]Q��]DAqAg�paDA6D�5!d_;kw'��m���������~/����w?�y��޺U���=�N�J����# ���Ma�4�)�Vk�'?*��L��+�q�?����t%�X9QP
�
E3nܸɓ'��?P�3՗�F��Q ,��ܼ|��@,�H�:���/�G��j��ɅL�inn��׿%ˉqA0�"��k���;�B���_b�7����L0�B��}F�ǌֹ���)�O��*�G!D�a�	R�<���\���v�UW]��x�؈����@�qc�����P��G��M���T~�E)֔����?�8�#A��������$��y/�T\L����P*b��tw'�`������?��l��}h�8�\�#�lk
rن��܄��=眷���<��m�-�G�V�Ga�'͛�}�z��-^�(�8�u��	�G��mӸ�_۰�-����kW��>9��*x���%�-1�4>��w��W]y%̏���+Yy,��*�JP0���_�$��.�=����F˜Jr��rΗ��B_z�@B �T�i~�E�r�T�B!�'<^�;�e�E����V�~�K_�mT���Vš�'Z�D@�  J�6m������
t��HA��C�<�o���f��+�$�-+����*n�]*kI@�M5�}����O����_�����k�-�M�F����2��#�ft����<s��W\q,u��W�9���vM �/f
�P��J�7:��#1���k��֮]��Ϛ3�3���}/֢T
t�V�9锓���wxd�c����zI�P�&���764̛;w�رcF������}{�lX��V7v�k�����&߲e�޽{�nB��w�SO=�?����F�����&�k�T FJ��x�u\�I4ι��k�����V�"�_L��,�T� )��g�+{����0B�F9��i�\E�/��b�3��!��4(�9��ĬZ�J2�dņ�.�j�$C�ϟ?3Ȗ���Pl*��P��z�s\+b��+�:��]�`��WbRq'�&3���~H�Q���[��4�]���>G��i"��ہ�f���Ml�}-�/�{`١^�H\)s/���' �¬<w���)v��1:F�O����n8ؠ	� �3"�a��.�*�����������$b�}��hz3[�tv�ŗG��/�ֺq-�&��4m�◗őYw-%[�l�2$���g ?����3���U �KO��e���|�#�z�a����ʉ�T�+}�� ���D=rPZ�d�t�s9���1��kp�W��ճ�:K�gd�e�c�9݆����~�̲Y	��R�� �$0��c�p��Ks�@h ��q�͉v��n`���>0�Y`˾��/3.�,�HS>�O`���ԧ-Z�_zt�,�t�ˉ�Of�C�!�R@)����/�U-A|)�)�'�pfz��~����<��
��������;-܁� (xro�^k+6�;�VX��Ş>��ݧc�����5�+����C�aKr,Jl�k����o�4�f�Ν��zk�Uv]Lr�8T	�&R+�7���П�|����D����� �]�jii����j��S��cL42�r D�@��C�Y^'d$z4���?�W��'?a���������}�r<~xv'���{���	ޡ��Cڔ�� �X(�� �g�С���y
���~H`L������_��KK^r�
��M�dh���4l��q'����s�@�f�߿�]�i��1Br���V�^=w�>^�k����w�f���"`�}��:��ӯ���a~J�*E ��[���7��<z�h�#Z�鷿���'ޚ�8N
�@t��i ��_�Q6�R�5sϞ=���o����YHU6�/��1dp&���_գ+٧��!�@�����T�}��?��1jH��%�(�*���G�Q�Ҩ�{6ǔz����͕3Ŝ(|������~ƌ�Z�G� 
`]@C<�"��AT� �C��{�G9���.�B��o@\Y��I��2�tꩧ�YX�6�{tO��x�vjeh|�O�Θn�U�6Wb��?�я�IxD]]=2Ş���!i>����J�wƙgB��M��%g�x�l��3%��f���-?�cD	zc�����Ӊ�Q&���+��r�qo-���b�Ig P@���_(������9���Ԁ@~mmm�������%!����g��^ReU��؞�E
[�o�t�S,A8-q��/nG��#t���g�)���:�(�-���ׯ�������Q)¸`�`���n���W�Z@p/�ń�M���{����dq[�!���I� >��#uV�HRj~p/�,�e"	Ց�����?���?���_~Y�h���M�ۿ��o���tC���,
^ �A��&��຿���?�=Oݢl>0i�?��]~�����믗���>�0�渖�ژ�?�я0�z+`�2_6�X
�ܭ$H������� ���뀪_�QzM>ٸq#�%4?�쳡�t��HلO�b(�@�!�~ah���]�n�ƴ^t�E��(h��Q�ߋn�'01s�=go1��
��1!�̫h$�|YP���&���P}������"_p��a�deWי�؊��l.��q��?���� + ��;.�z����}�d+�H�\���|̚5��C���q���R��`�0A��LN���ó�|9|	��Uu&�c޼y� /w�P��l���'�kf���n���e�ᱮ=�!��i�bS�>E:��R�����&?��P��~������_��\aC/ �z�����o~��7��(esu�9R$�[O�A���a��y�e��cr!���;�+_�
�n)�]R��h�f0�pB�Y ��AL�� ������f�0%D�+�8;����s�=wժU`kn��?����
���7	+Ҿ�����>���+WrI+vJ�T_s���|��+�łb[��/��p�ȫ���v�ZU�a���l&/�0S��f���;ȏJb
R1��656�~�i�׮���nۮK|h;1�S?Vq��Z�vu}��ߛ|�[W�}����Qow��}��t�1��j_Ͼ!�t����䷞r�>�ƿ>�m��if���Ɔ�Ãeau��8���&@ѭ]��O��Me�*T�
RZf��cQ��� ��>;z�UW~c��W�/_^�j&˟?=��S�B��j��@���kπ.!5��SH�f��gߩ�ft�"�G�<b�e#1�j�+T4��s���,]��.K0��B���?���.���/+o�����V-�O@m�:�*'p+�A�b��yt�M�@
<E��d���']�B�g��n�X�B�d����3�<�X��&�Q�� q���ǘ.A�^I͂`����?�D�Hg��������F\�h��߮�W:��)EŨ{~i���t���M�:�S��̬ٳ����N�H������,x
�cͦu����#�~�Y�-�뮻�:��li4x�eƌ�h�\�Ƿm۶~�&����U���a&��{	��4f��5����0�
�38%w*�D87��+�<x02� m�Wx�|!_�|��^z	Tr���߿�]���� N�/*ye0����'�|2�����e��ٖ��p�9�$o�l��/�{������;��\��Nl�*�	�! ��g�Y9�_Ȩ7/��ߔv���ہ5kE��>�t�9���b�`fwo��ܛ�:s�1�^z)D��ŵڧC��E|reщ�Y���4�x���o��	ɋ��7?@��mp��@�|2���z�2e
<4i�_�T�#cQtX����t~���[��o�~2x�#�����a���8��;�=,ؔ6t�e��l߮��654�zz�<�.�b�#��^S�&L��W�:�yP�P��n|:�)��T� �K�=����޽���ur�AL��(��2���Ϙ�/~�Г�1�.tl�ްe�y�8A<�����ʒD	�_�l�Y-%��T��M�4	��|)�TN�� Ј�`L1��a��ѠyN�%W�O:�$�t!��� Z��-��q���o}�[���*�tnF�ե� h�L9�<��}d!������ŋ���c�_��e��.�䐓J�*3�����,�s0��ui��e�D=`c�Z�v�;��cQv�s9l�!i��掎���0X��5�x	o�=�^v,�����_("���&À�����=�쳮�"h��O��w��1Ne��p�K*.�[�7װN��}�Cb?%�"�
e���r P���w�/�P�GO0�c�=��L$q|�(���/��/�?�8���^\�j'N�$�e�(0�%B+p��_{���.1�7�R_r�%��ܻ몑��1�>�o7v��/�߹s�h.��(��YR���s��]Y���O~��{�L6�_�߾^�ufx���_��pHB��-S�Nݴb�U���=--w�y���K?�A�l�+�t�c�f��q>�������r>�w��|�B��J$,��䃘�뮆uCݞI{U֙�d]p�O<�Mlss	�$��LM�A	��(A������?�M7�$��ܒ�ʮ��~��9R}+	*�[�c!�[�1�"]�~/��ts�2GH"O4��IKK��_̭�� z� t�A�	�g�}����%���#��S�����/�V�Ǐ��O~N���C��^�Nh��8��4����pm��@�̘1}`��C�%���hpX���裏
��|b	*
���r�lL�o�J)�l��f]?u(��9�h�}��=�PWw�iӦ�M���V�M���qUFGz2�4�/,ą)!C:,-
��@r�� ����Iߢ��3ԥ��ަo�f�o1�Q�����9�����U$*�N�B�<j�( Q�rҷ[~�γg���m��x�����-�Q��a8�/�}�{��s�ɐ�&�������V�*��8���|�ĸ������6��!���i ������E]��$�(��$�^���{��:�a�]eN�)�g��!p6�s��Њ,>��;���UC�]����
�{]J�5~�>}:p3����6���U]��O%���0�������^��<��
�����m���\���w�zSgg'���?̺[z��uz�~T�7`�,�"�{�l7���K�G�$��_�Z"����pdM��vG"P�ͷ�)9�2C��+�i�JP������ѳ�g'RvɋPD>��՟�R�� �ϙ3G9����^���h��j_s�5l\يyºl���8��F=��/��ʊ����!���|��܌Z����?AB��R!Az���@��iA�f��{QM���h	I�k�-��9���ɓ'Ã�}���
V	'���͛7�n����a�H�Ǣ�A���&b@:��s�ެ��� �V,G�}V��a���Dj��Ig�vf��m�H}=W�Dbs6�|�5k�r�:ٴ�rȹ�+�ZZ���aK�| ��ȵ�������}�рbƪU�|��"�lnn�g���}e��:�,���f��m�Y�Ï@�*��S�X��*�A����/Q߮��Q�y�y���% {|�	`R�7���w�Vt�{����v�;��Κ�;�]�>���/�������^�з��<̙>�mok;jo�tx5��|)�y����Q��)���sws����m�d�l��F���7����M�9,h�3yА��v�ޫ�:7.xN��j<���=q}�K��o𳾮��3�'��h��&y�OP{ي���.�9���T�t1��N��Ue����J̶r����R��3g�<���i8ݸ���D�(�����{/A��BD��%�H�]@Y{��t�V^6l����t.�&�	���%Z���){%p����&�t�}f���"�N
)\�J�zᰅ��z�k��V+��d}`��l����S6J͖1R��|��ɚodO���F����̉'f�d֡3�8㌛o��V�7�=��h���&L�<y"�?��X\"��xvh�����(��7w1ą1��y�Ə^��m׮�[�Å����S߬Û���"�8dȠ3�8�PY���R1��'�x"��n����Z���) $��\\9"��v_5T+`�T��a$��/���&�4���Ip2{p{`K��V6�,qc
G�w稲�\Lu/�#� �?��#�Sɍv3�������-|�Ԝ@��3P/rC5vfB\�#�Ẉ����Mt��_A��u�|B�
�H= =���SO��o��յh�`8Sh �� �E6ܾ?P"�& 8Lh�0=���Ag~��#G�x���,�����z�)�456u�t���$�����oX�DĺPu*��-��s��R(�ys�`��T�0i�k��	|�v6TB��6}���彍MY4�;���:�fzR201F�,���۷{vo^��'�zL�O^��3$��0�� pZ��b[֓�������K�<��*:�ണ�:��GUN9��)��ѷ���Ċ�c[�%�Ô�t;��D����0*�Zj�WRߞC�چj�E������/��:e�ݔ�G�k�\{h�r���W����LYr�H��+����u���B�.�Aڞ5&������&� ҡ�$֋�p[MT�����U�M)����A2�ʊnU\nPA&`Ĉpn6m�$�?\8��$l3l�g�U�K)R�����m�6�y��g�1p��]�꼲~p`���Sl?�0<����8/&��%�O ��ڐL u9~�x��Fe������ࠉ$�zft�)FD���W�h��&�)��>��ג���&N�x����T��4z�����^1�q�@�0�0mv <b�m&B�����E)H#\�:^�s�����V�jk۫����Z	��C=N��~y*�A>kY���K|0���"�(�8c��e��
�{1���-q��6GČ���W����|=�^�8�S8H�$@6梎񒀴�J�#M����{F���~���c�%� 0������{3���a!(����b�\���u��IJF����N�q�u�G	�޺u�P��*���F�+������'ɐ�C ����nӵ�50zf���3�e��cƌ��߳g���M�5��z�����w�K0�r���˖-E;���*T���c?ʏ;Q|MF8~���#���!��2_ &o~�DEI�v]���P�e#��wvT\�]xA7�2\  �Ȟe!�r}�
ߌ5]"�j���ng�0�&󨾛���ӦMswj�۠�E�jP�����bj����N�x��]U)�Z}�m�<z�B�
��[@7n� ����~���(&��:��f������%S�E��8��;�s�޽��VP�z�;w��V��]��E���J�V\�h���7T��H�9�4jp�1�0R
T`�"�4'<���z�;8w�m�mݾͤ�UP�=�b�<=�;���Im���ښ8;[�2@'�=�X��j��*={t#��l�l�i�5|� ����۠������,����IR���ӧ�mD�ju�Z��+��^{��pĶp-=m�;W�V�_�$]��)���-[���h�\v�U�r�]b�y�邏N���[��+7��@�� ����/q$D��$�dɒ��ri����{㞆NO墖�_Zl��#L��/2<Ӭ��8�#_ru4��ye��Ȥ���}(HV����r�-�ڳ1i�?1�_���^2����B��
�-��[��Mb�^xpvu�����-_�����S �|��R9�!!PƉ�d*�Z2)�a i�=��4H�_�"t"�7���l��H�k�3u�3�K��3	t�%�I�)��5v̖m���Saf��Qsg��G�L��l0v�� ��6��77��X�:�sy?WT��� �G��Y2t��@s��kJţ�������<�l׫�r==i}��a�8J���Zƶ4������T!��M�m�Eh�d����|l<h��C��N����������%�&��k]{�U7�|3�p͕��	0D�X�_�
�llAe����[�w[�5�W��a��'}���W���I��Gj��x0�n��Rq��B�+'Ѽ"Zq�,@��v����&�:��<$YpQQl�r45�i"�c5qd������	&�%��,�{A��@%�u�с�Mp�'�ߵoȒ2�+�k5z�u��(	�͹S%|G��n߃�0u�de�z{z��9�f]�K��l�@a]!����AK��)�����(p�M7��Zx����<'K��i�
`br-X���U�����d��b��x��}{��^�3ˀ_�wg\x����\��-�@�Zd�`�����h��p;Ջ�7�\�� zn_���h�\�3��fT�g��y�)'}p��R�ZZ0�o�`+G�������P�rł��,YX��˗/�u�6����:uŤb�2�-A����5�i
xYy9|؋//�hߛ���-W�-^�b���A���/P�������S�T_��av����'���Kg�=,��z,�{�: ����Ÿ��y�c��T�`]��O�w�}�����۫[���b����>�9��0�,4�/��W�B 8Af��)�����lȿZ�U<�ۓ��	����KHqA�K����X3SgI�����Ud�B�&`�SW�@�r��Y}�l�N4E�X�bu��;E��hs��"�&ؔݮ.��^��,�f�V~Y�K40{^!�6m�6�2�u�w}�$&�C��}�ᑸ~�8ل Z�N�ʮ,�41�_�:0�R!Ԗ��� �㤿�/����M1dsȹ��X��ڭkI���?��s>O�HΦ=��{Ɲ�2�f��
T6̦�^jc�lK�����ݭ=��vխN��
��@V}E��=���P�m@��l��s6�q��j���o�L�8�b�i#�8�pϼ���a�"e�d�}�6_hX&��#ʲ��(�SX3>�ł�H��]浄NY=�F�H�Z�I�g�<Y��Q6��n ���q}-҇�+�2�[��V��ˁ_BY�+x���ב�Bb�� p�o�i�Wř�2a��?f:�W^F�Pn�0Eng�~Gz%�X�!�x�X�cJM���;+TS41��<�\
H��Kf��^�k�{�R�pg�U�+���C{b��H ��a�����i�[�.�gչz��eɇZ�$����W�؅s��\j�+�<������W4<�J�շۣk�v��������K��y����x@��8����ȯ� L�K9ի�@�f+W9聻��q��BA;�L�Z�j���:;;��޾��8['�\����ď#���rT�𛮝M� �	��S��y�xh6���N0���x�.�7)A�h���.���;�h����Ĳ�Ui�ճ�0��+[f�n��}'���_��T#��EƥW<���Fۇ����Y������H!ct��-�"��� L"����Bؾ�D
bB�19�V�A�.���K�z�H�8�Q�g�Q�0���|�$�E��z�%S�f;�2kdZ�%adJq{f$�����
2��mY�G����p `QqE�x#�B��X+�p�+q�/�{y�Iu�G�V4^�H���{�mJk�=�Z�'vM�߀�G�Ҥ�͜�f
#������/��Xg +��
f	�`B�$]^��&~!�ZF�:|XOo/|�ǟx�g���;������ՅH��BH���hI���b80���θXLw4��0�I���Ž[�ޡ����Rd|!U���֚��v/�Hbп�Y��TU&Ѱq��s��,}&���U��; _պb{տ��L�Ua;�r����s�eu��gu���9-����k�΃��*�dy��I�
�=��&q��Zp���!ZaJ']� i�t*LO�:-��gR._�ԤF�b?J	���%�Ї���rrj���c{ڃ�  ��Ϥ}ʺ�4֑���	���0ʺ�f�+h�,��8�_���S��y��½�����/���V�j�L�C��z����)�{����i~�G����f��W�l��ā���$w&�(a���D��?qR�%Q���/_�\�E�t�}��Jˉ�M����^�w=�"�P��>�t�LF{R���
M m�Rp��F&e�=+�R��n���=�V�h	LL���w��4��}P�ֺ*���F�>{'��b����q�^ʑSq�� V�+W}��ܡ��se��y�ս����xy� �� ���$?{�$�����I��EM�O����m��;';<{���͛��2�����B�x�Ob7��	n�H�$D�����w���1�}���===�w��R��׾}����X z�,˥��{{E�$tDk��w���&U�����V�FC����nV�r}�(*��v��[;�Ƥ�N��)��O��-�ٳ���.3P���,|���M(Q�|Qe
tt$	�u:���3Y�VX�MFV3�5��mݺuР��{�u�zWg����B��nmٲ�����:���ޞ:|"�ط��0��7�Z���6mb�@������;��׃ x��i3MTN�����ݽT�A7TI������	øA~��-#����ʚFd�_��W'��|z�E�ĩ������ʑD�<)��u�UreS��箮�����)phR� �~;_(Sa
݆4q�#F�hnn&{�
-z���7�zH�3q�Xv#*%�ٸ�-}��]�vIn��h��j*��]՗��E�R�*G���6E6�(|g�/'��}H4fG��J���8F�8�I�y������ջ˄�od�����"y��Xy�~�
ɺx�����?1)^��*W��~�T���ڻ�り`&���V:DdO�́��S�WB�z�v�򌜃k��jU�]�u�ǳz� �J2�̌3�l�W��@���~�z����k@Ӏ�C�v���tI'�{��y�z��E0S�zj�K�l߳���ʂ'���8;��5��@HL���+Q��7�m܈����w�<{��ETCv ���o�B�<��w
-�Ԡ�xu}cT�3�!��qR�!���܀B����Dw��J��i��W��M�0�>�B�, �����n��0�e ^�B({+�V�4l�'�G��K����$���5�� �S������uH�������o��S8i�x�2PoaE؝$��?��S��tg"6��=���0r�5��������D��
�%<���,Dݷ��2�: ��쫯�
=+C���`�ڵ@���vV�q�n��[�p�_䥞=�r�ҥ�lbz����U��<�f͚Į	�Q)(3U�n}��|ى'����}�b�f盔��$�S?�C���ثJ�b���{������5�����Š��ޓ�ѪΝ�[�N:�Q�͆M�l))m��LiW��l�RL�j�&�T�pSF�{r�׬��ӡ�3(�V)��u��^|(F��l*�~G�Ύ=��R�1�����yU��U{=`�W^y��\�u���>w�N�޽{��[��E���/�ґ�ئ\ :���Z��L{�����j����-���k�V�eܽ���dݺu.��m�3�Z�C�����Eav�?ǣ�E����^�Zaw=6'X�u�Y\�Wu�whhsٲeг��6q�@|����SԠ�`l��I���u����c�������*�y��T�n��}{��t���������<6�S��s���,�J��ñ٫Oy�������<��2s�^�Оz�`,X@P�*aW����ː>80.2P5������@^y�-*)�Pt��vZų��½�]W�Zá��Owt�+t;�0Ru�������O"�;��x�]v����@p9v����`�3�8�꥾IP���2��ֺ|�r��ٳgW�\��"b�;*�O�S	�sGxݘ��Ln��=X����:{���TQ!�|�4\�B�4p�.p�[��Bgbs��	�n?tHp����4k��l*s�]�֎M*H���d�{��{�g���W�c��^z�%hi_&����āng#�*�E����WDQ$iW�];>In���8?���p�<[���
s�2���x6�#�'�Q#G��ύ.��sP���T�b����ᆍ^_������ݴiS����]�v�i��Y�ڗ5�M4^���>��\���~��?�4j��Bߩ���U�p�(��7�ca�G�q��<��y�q��B�l�g�a\`h��a��MFT���E���0��}qb�E �����{������"��I�'?���D�l֑G)��Ef��&�ӟh*r��-�joذ&S*��hɻ\N��zL`C6	(�E���>�����y$Yb:�T���&���D�7qB��c�0}��ގ���,���~�.A�6�hF:'vv��ؔ>ķ���n-��f������S:[�TN4�������r{;��)�/FEe�G:�$A 7�j(W��Ihe�96��gŊ��E�+s�!@aII��I���A�ds)��Y��.Y���u�5���o�d1
������}���������~/�f~�~p%
-�6++_ʲ!@00���������~ҷ#Tǟ���:�wB�ð�~����݆(A]\^}���<�ǍԙG�&�S/�xa�J_��_a��k���N	�*��K����n޲��4%��T��޾r��2���@x�s�	�岤h*m���]aJVJ����)(�4�Cn�\P�nt��3�b5e�`%f�V�*�O��'���0�Yn�m<a÷���8�ۦ;��-C&6VG>OlLG=��O��=��v�Z�U_h
��u�fq94�2�����mne�j�����$������5ٳ�V"{� �sĒV%{�J�ȧ�8!Zş*��n�a^n�q��`5|��TsVq���x�_�Të�x�n��,!P�rtP/`B�CRʐ���73U(�j��d�}Mp,a8��iY'�M�����{�q��4>��N�zPScS>o��Jy�)��4D�=���6(�/�8U���m!��g�<��pO��t��zAH����A�z��*� QG�v�vp�h����NbCh���+p�����g�s��'�Ϫ� :��E��g�ˌ�+Z�%�:�I���U�oݺ�Wm f�Dk�?�<���X�}v��.Ђ�b6
՝t^ޅ����%x�q�*t��e��<��ÐA�3�^`�'M�$��:��dO)F��Q�}����P��-E]�s.4E
�z�J']���^:6�/�N�2��� �	����Ħn���F�P��ܳc�m7�|��C�L�X���d���Kn O�r�I�I���除 ��?��<t��D�&��/�Zg������o��� ]�B葧�~���$��a�����u��=���S���Q^�:pꩧ���kd��;12j4�����M!������F���;�8��
���~�/�9�6J���8����.L��|I�DI�����?m����'�lVs��U֏2��;_*F;_Z���E�y�U���{�c4��-1H��9?hi�ջ��|��tWC�}��,U��Lz��=�E/�il2a��/-)؝�~vـ$�m����C�]�il��t6=6��Xg�;������J������}��G�|^�jB����s�(f��ׂW���{ϟO=�8].l�ߏ-��Ί�	�&��82��/�uǝ�[�i�c<��3��2Ǌ�ҤA�n��V�B�Hlt���I����+���3KA����
@�����_�����3%���)��ٝ=� ��7���ˊ�B��.�3w���YJ���r�q�F��Z�\E�@	��<���a{ܤ�~?��h�裏B ��V�Fw�M7I-Ax�]��!�|�Ͱ (�@z��k�<�L*P�k����Qx�|'G������1�]<2eQ&������Ϟy�ݽ���,��Ά�� l�:�==�%s�D�&������N5d������C� �Nh2l8� �={���ׇN>�̬_,E�|�汴���ā�����C���-���~#�741ܫ��k-B�&����{�;��w(J���\��x�^;�yꩧ`���|W�q(:���?�y9��eo��K1A��7�x#�'��܅ Y�����u�gH�KbS"�W��K�_T0��2$7c���v4�ĉ�Y����(�9D۠	 ,���p윺�~�wΘ1����;M�Y��g���׿�e�jVWF}��B=��딜#Ô��|svO;�:�����`�!G�z(#��8�SKMzE�M�����\ӤX�`t����H��i�ԩ.���SN8��e�>P󮢞��K�To��1� w߾NP��� ۝wݾ�us���u���}����2�Ò^	V~�'���2e�ʕ�O8ᤜ��2���RS�F!6��|���i���m���׮a��tx�7�p�W
ĔZ�.e���0��`K��)�Op;�.40�+ ��:)�̂�h_�ݠ����~��N�<مC�=R]9K��������x�x��	�%�nRIַ	�vNJ��$�'��8�1x,0y^x!��-m'% G��?� ~�
��/a\@�3gB�
�*��"�Ch,���򗿸�������e�z9r�oإej<g�fd���cպ��7����$��7g����~�ʊI�bc*z��kDz�,�L�y���cS��8ڰU@�����e)b@�s��e��0�������a����͛��]���#�����:��I���#]�0�x�@?۷��Q}�"�+|%��͕�_����r�e�]F!w7�v����!�0��w��я~T4o���8�N?�t]4 �&��gi����i.��'����
�w�I��^c���޸!��Ky�͎?~ְQPĭ;Z���9~<�T*ݥ�]]�U�Tnb��[� �N��C���hѢ5k֠׍��Cy��#?�YZںD ���t��G�C���
"����2DA��t�TgM�?��%����о�=��*\81�����0�����^gN�g��c,Xp�����<|�E�P�	g2��S͹�w����;a����О��e���p�Eh
&W0!^�qbOg��޽{AɃ:h�����5�&A����Np����z�8�+� �|�������qu��Wx�$�z(ҤV��3{��g�x≞]3��M�okSW�A ��~�#������f͚lJ4�r=�V������_����N���2jԨ	&�c�W��W���׿��2���%�T�P�5��R���3U�@�F�W���}�{m�w�V �c֡��Ч�;w�#�<�L�2�*���Co�Vv�$a����mH7�JL��U�%e40^��KHXW�%v�<2��+���w�b��m�����2�5Uh5�����ubs�.���M�U}O/"�# ��?^x����ʣ2�����A�����,pח��%��ok���1Eel�����_�M�#}P�@����� E�XJNUviEB��g�y�W�L���� ?����ϟ?i�$"��:��c�=Y(��V�p?t;z��o~�g��Q��fhBB	�
��34��4ެW�Q�ke�����!#S'M���������E�TOoOcCc`b3pO�91�9=ݤyf! s�ha3˰&�}�j*�-������A�GuԠA�0�x�;���=���wVh#���A2����9z�;�9g��T�!�G�>��6D�����,��ٖ���q?�#ƎK֒�� 6B�ϛ`�7]eϮ���V�!qx�3��K����_�UȘY�)t�g���<��L�>8^婧�������l��5�(S^�	V��{���2[D:�"f\Ry���=�XhcWe��؀:K�	9����V��%{���'?�	�N��2)���s�%lh"��ڧ1������&#8^���t�ww�fҰ5h���M/��FL��m�7�6��dw�C�$[����0rI.���P5K9����xA��a:�ﹱ�������}�/n��cǝ{�9h���e�o�	t����/�|�l�$��:�D��׾�����)G/+�e�p�0%P��Y��ei�P�a:t(H��ge1�hF9��O���&V��ꫯ��y���������$Q.҇��Z[[�7��n'Ů*�?��P���wƌs��{I�t�L>�[�
��F�6�%]V`�q�>������6�}����C�r̚w��ؘ��O?�����~ԣ��������[���6DH������i[xϋ/,�w���J5��%�����-�v2dM���Nlڴ�1�4�a@��ڠyܜS�ف�.ذ�%3(�T�7����»����o��_!�_,1��=�����1�0�����幑�@�]q�0�s͕E �yw�څ�jii9�S�WT��j���#�����}�d 2����b�&���F�� �n��o�y�J�.\��?�)s��.^	����+����_n6l��u�ب��V����gp;zR�,�,��o}�[P��z׻�Ӫq"���&J�Ca��e�mE���!f�k�9r$�Rb6q�Q��� �	��j��FCq?=n�ꪫ ��>j����i��#�A���P�O#6;�cB%p���G C�ŵ�6�r���t��s/� ���ܜh}�Ż�������"��<Q��{� �)3�^��Xȭ^��y��t&�8��o���'�(?a�Dx0ɞ]M�M1>btҟ���T9p��R'���ab1S��X��IR�ĺ��@�/~�W��̄j���̺u뮼�J-�0yb|ar>B����r#��ѳ��\�@ӧO���KA7	���u��0g.�F��	 ��p��=أ~���Ĵ�ٝ� �����~=���)'ʞ��+q3^����3g������ImY���̇�硂�%������?��q�T��C�/�f�����3%7W_l~�A���s��*��ʕ�Ya����rD���t:�-�q�}�ه��ֶ� ��2��3�ll��zt�Ӝ��J녅�)�m���˗��-�2�W���+W�f
�|g:������;5t�~P	�<�3RR��/G�y�����<�N��Z���W�
p=�/���-A̍�<��s�04W\ �K�'O��'?	�N�0x��~B4�K���K���٦l���C�0�@2��
�)W�rĦ0��L��H�����/J�c֬Y�e1!v��J0�^{-s�gML©���x�嗿���c� Js��p�2���1`\!��S�fV�q�S�N���7	�F}3�g?1��v�WbRQ�s�8���裏���G�/�T�(_ȦS;v�_��ֲ��u�)�����t���G�Jg����`��A�����'���R����e�eU��̧�=���C?\�t)��S6)g��$�`v��aqE�T"�5���}�Qhp��!�M**^b�D0`> �,�r�����q֯��:0����Br���S��󇷐���~��2 +C����Ϩ��rD�PO��Iƽ��ܤ�P%w�+����w t ]J�6*ԥ�Ju]&�`�p����_|%��Y;<��[�9���kVk�h{��;`{N��}Z���ܦTSҘ��ttw�\:gq��]۷��E���^�%�T��ݶ/=�����_�����p��۶m��s9���G�A��mR�k��q��7���;��8^a3�4QF��:lch��ܴP�;�9 ���P��6�8u �4ngGYt"�{�v8$w�uW���xHt435��0�_��W�:�(����8(|�[p�< ��^S����pGY�/����`! ��3���i�|�ۿ������Ce����	x��sυ5�:�r/p�4 `k�ԉ�sO=��S_�җ M<�]HۜZ�k�<����Qz��x~��_5jc��개FɈ,Ն�]������g��4�����R������|���LpA˸r���Dw~ӦM�-����5P	�	S��	�\�+�t�.�T*B�`��9� $v�� 7��
8W/Ad0!�G#�+��ך\މY��E�x��˗Ȝ�r�����?d�2q�e�&��D�.��"#��Kl�r>�����E|���SuW�����/ql��HPR��j ��Aa�0��Q����4�(��]`R�o�a8c`I=Ml������+����:��&Vzs��49�c��#0�/��f�*��a~��#&�"�@;��7�t�w�R�*I.� <|�=�@���L�j_��u�!<"x��=�R<LѐO��n�A�)���`�J�1�f�N���6����O;�l=��L!��ҥ��k,��Ƌ�yf!�����	���텁�\Ç9l����,X�n�H1:v�i��t�折.dp�ƍ@�O?�4�������r��S6g�FE%3D����<�BG=ƀi-�K??!�x��.�̲�����|n�!hkk��Ռ�u>��������t�������p?h�bB��Kb�NVM ��i��r����}3�i�{�1�d,���#�q��J����ߠq)H!�A��(��?�	�+�/��5�����Ǹ_TR]$f���2���T���&*�R^~��@ԧ�~��0"���ƾ�/�_��4@��Gˈݠ��MkN�qj���]�{�n�"�m5o�śBR^ռ�>9�!���-E�������%}���2�.uEPxIT�<�����GF�eg�8(ʄK1y`.3���U\%�@#��;w�y>���Ǎ;G\m߾���7�1ln���rӿ0��`YL�[���oȒ
9�������o�T���N��>�!f�IL���m�a��]�_m��~ �~�a��%��+��5���J)]n_�a���ǛA�m�wH�{1^ �����F�Ͼ��g��	�Mlj�K�)�_l3bLז�/xj�����M=�(�7�z2��; �V�mY����gM9��RSX|�֛�2��Ӿㅅ����F�����,[V�k�^����??�KV~��<��:��`��Q͠�v���?��C		�b.�J��>7d�啘x��Xb�I���8�&Vªoϔ�,|�?; ��9���?TGE�Yc�7e������0+��W̃��6;�7���z݃Bd�fX%v���9�V�#K��T����uދ/���ڊxN"1Э���{�U�էO��L!���w= ׂ'j�N2��={�{�9�o�� F-!#�4�����@�@�p-�jc{L�2��} kmme�N�\�Wڂ��CC�ړN:����}b1��?��Ͽ��;w���`
�g��tw��߰	X_�?q�k�v��7>�S0�CZ�7dR�y=��t�cgۀƆEϿ�����-��`ks�*�����ʒ�w��9�<���p��]�N,օ^&�""������������`��/����@}��*���?�IQV��5�s
��%e���G��-=�3��!L�+���3xR��LaS���o�m 7���ի?�Oy�<62���`�?��u�]�a�ǫ����z�|�r�J����׿���0a��].���0 �a�L���«0Ix�3��`"�t���\�c��2P�N������3y�x��0#��~;�Hn�|q�����C �POr5��A@@��Ì�P@H�/_����BL��h�S��ޑ�Z[��n�,�ip��7=��c�_�*�S����ҢO�I:��C4^\��S,p��򊆶I)?�`7���b/*�u�t.����F�G�f \r�%�Y�n�.Hă>��W&���.�Ї0< �����w�C�i.�<n�,CI�v�m�\s�C�ID��2��s���~N#z%�����?��0`ϫ%@7[�٘|�9��+���2p-(�2g��a��J/�8)�b�h
��G>��O�e(n�c��	��*`����a!�� =Q6Þ��{Ŋ�� 8�ɽ�:��wB� ��x���̣ok�"���E]����ĵx�b�	cN�&Iп�I��!D�	i ^ʦ ���{�WӺsG�����Ѿ&�Q��lA��D��У8p`�ġ=��2ʛ���Ţ�"�Ӳ��_�<&ISA�������@�����6`�ѣG�u�*`P����I���K@
�@�j.0!�@�j�bF��DY�]`���{ ��w�̙3�me<{hX�48^$ֱg�N!����}t��ȑ#\�'��'@
x�P%���!�Ӿ�`����<�3@�I��U撇ޮX���qْ��^0B�X��.	���\���L��3q�\t���[�|Sӛ�8r�`��m���	#t ����k����rx�op���Ӕ�\`^�����t�#�iÆ���Uڟ��g=��	'�0{�,���C������
nF�A
�bE�P율1`�-���w�c�!����\�5�T`�%K����U�Z*U�+�EM����.�=�/$�BXf�F�;��a$�(b�A.��F��ɯ��c�=�֗q>�0$`"~����I��]�RL�@�P�hv���`x�8!���'�x�3�	�{k~�}Ð��0���?��Aq��Y6�nC�B�!e�G��`Gv���[nd�5jl'�
�n��A��N= u-i�%��� BB�mx��g��$M ��h�r�=��<nb��0i�H�B`	4��K/��kր&-�G�{cF�A��ѷ��W=���m>���)��q�hdoW�N�O��v��|?��طg/�(H�U,�[8�G����t��s<m��-K ��9���/�	�'�a����|�ɳf�1b�4�߾};�ؓO>)�[�S���Y�s�t�_�UV$�3g fˀg��g�}d䊊���˥���_e��P��Y4��π��K�6f=g�_�)s���%^�Q��h���$�|�f��)��K[KT�P��Ba.�k}���cPb`x4���\`H�_ƃٙ�&�R��c0Y�N�- z�3��'h��c�=�a���W&h��4��&��<n�����8z���MA;;w�D�0�RAE��W.]mc����KWa����!�R�.A�S������Ŝvqs&��a�z̦�L�t�^4��׼7�РO��Cg@�)��z���n���g�!'M�=Fnǻ n�|��:�����^�����P�x#h�B�ar!\��:��0A��p�
��ؠZ޺u+f��M�U}�z���V�6��=! ��~�3�v�U�����%����@Fn��t�ke��nxô���x�Gu5 G�A�a��W����[�I��dKr�A�#.�@a8��!gϞ�Q@4�P�#�/� �ʍ�U\⢳焎�v�	�/�Z��� 8�A[rьa�Z�ȁp�gJ��k�E�� � �tu Њ�O?��Nm2ܞml�h'_翕5���h����z�/�O9^���&I^[�l)����<�l٪O�^?b�.Θ���z��/<�?S��3U�Ͷ�R9E��.���x�[�9�6C�d,�:j�س�<�{eV	�ܡ�� �,,��g�DET��%�be�O<��0^�h���CtU�uָ�²-Q��s��gS��C��*�'���I��I��:��7vL7W����GI�5NQ�X��Z���ڤi�|��Nm�SZ t����Lȹ�w;�Ls�g����4~ҜZպ6<d�ȱ#Þ\p�D����{��4�!`�Wz;��e^ �`q�q�1�%��`�����v���אd��:���j*�џm��7d��v�+Z�i�_4�s��/�{���_�y���ց� fSV�fOW����8�,dW��EZ8�$ ��١��P�EN�qX1�G�0VG�z6����D�%��AY�(�B�?��yDL� C��P��/�$�S��YH8|f�jg~��5L/�UBɬ�(��\�+����l<| �:��r�c*�,�.���/�W&��i�V������)MĎLJv�� Rk
���n\�IL9x>�6Z&%�2;�U׊i��"Ӂ���������aV��%��S:��LX��²�����	����+�W̜9*
���_*f��5����Y�X׵�:qls璨�Kd1V�>&������h89�6m�vΐEg c��	��7ވ���E�y01	�ZO�������0 !Kl
�`8�v���a�`H�h�#�_����\��2*]kFI�*�d��BSh�	 �ٔ��ؖq[.����'y��s�=w�q`�gK�	�`����K �Q}��M�{@�
9b!	�46E���^������\��̅v���8x�����fUw�;0U�(M2@�����vh�����Y��.�XU��E[��H�[o�<�(�6���N��FH��:_ӜΆ�|h���Ӡ����f�>T��L�a��X_��s�\a��3�m(8�/��p�-o~�رc�y>���q��A
���[���pJI���εkV%f#^G�3�L�^U�s�d�|�5U�Kp�pN#�l�r����P��L(	*�A>E������h�$�j w�w�}�����Pb`ڣ�oḤ�GY�En'��	�B�կ~�-�MF�c{>�[�L9��JUg{�2��mEP�Pe������čbpȢ�
�L����z������T�+zΘ���T�J5��V�^p뭷�۹�@K��	�F���F+�bG��aL�C�)Tׂ3K|��	L�Δ�s=�Tyf#�%�dOgONy��T�����d�_�����tA�C��Z��r4���AN���]�k��U��K̖|e�a����k�jj%�,V_�K��&zRQ��<!�XR����T]��rs�$�Kp�dv��q7B&S"Э��)Ñ4xb$�2:�B��ܾ�RpŔ��K�p�R��3��U�H2TyG��&���M�Yc٬�/�%�� �q��ɤ�Ҡ	:�=�!C|�����tt��x�q�GL��5k�3O=�Q 2>�v(��L����j�Z��;v�ھp��+*� {UW����vB;�F����2���We�0�g]__�ء�~ϖI�n���q ��B�_cÍ\�#]��S	�-$ˁg�.�o��%̆���n��5�	���C�痀/�ز����'2��U�E€#��C�Ia�W�JTg`vq��e���>�Ј�����dԀ��b!Z�	�������&}�\d�NT�^�-H����"W:���Q��B��>��ּ�a��)��2�F����0l	r�x�ĉ�	a����Z�q��R��y��g3f��OL�)S�t1�H�( �Cx!_��v�;:���+��.s	��ZzN��B���{|��R��y��݀�)�tF�@MJ��ll�߉ ;RL<S�HY��l,q�Wz��6��)DYT6陝��EVI�-�`��(E��%�FB`�s�y\:�O��w�O�R@XdA̢��$c�+o�SG��l�U���"d��̔`>��ّwպHJ�եu��������]�؅v/_YN��>p?���`�95���G�/�+V��̙3y(Ǵi�d#rT,�fH%uQ�+̝;� O�0A���Q���X}[�h��W��!me�L(���_����Z��[�Y���)���%���L���"���Ll.��:$�oﲁ�TQ6
#K�,ں�P��z;�� V��+w�UŝH�)C��m�i��\��"1/���� �?�:"�}[�B\�g_��Q<Wx�QA<cXY�+fEYDW�'���ca��v��={,L��W��p@��1���'NO>T�;~�� �<h'�u��=#;���&�6���ܵo����Z)녲��P������EgM�wv;)[G9��нD��Vwq/�]���/}�7�[�TΊ��P%�P�/t_!�%2s]+%-�GmҤcS0���\e��J�42�,�H!W4Rg���GT����|S�1b�G���;��>���lcw�����Y��p~ʔ�3{�:�bGP��6M��:lǛ���~��k�F�� �7Ν���:�x.eG�/t�l[���m�ж'j($��{��U�}Ş�Y�:������ٝ���y,���/�q6s��-rL>)��<��| Jcbwh��;�<�$vd�v�1r���-�n��p���)��)�
�:QxX��`��2�kk���U(e�>����{�=�Ț�E��<�-��@�.^���RPF̉lN��@�%�����R�Rמ�n_��%w��̦@�>�~������(����\>@�j)*�G1�y�$��'��ի_�O����]�f-�h׶���v�Qp�s�����ooG�P*�9��躊����81Rq������eۙ8�\�'�Vp�{�x�����G�D��B�V�UN�8/�_�ӝ��ߓ�V�մ�p�[mA�e'7��B3��`�P��*��3[0U_"�W�"�EaW��J�r)��7�H�^�7�ɥ��B�(
�:.Qe�-(�����Zpm̝����)����Ty}Cy�ʞ�
t� �BA���^[9i�T@����)�xi�"�h�җ��=������A��v��~C���HoJ�3Q�t��֭��Ϙ�����f'*�3�m�`[��N}bj�ŋi�\�tYȥ��'�vJDRb4.��P�5��ɾ��T��ޮŖn*�
�W�w�Y4O�w����݁���D�̊2�����k)T_�t�W�9�������S�r
u��f��q��±��.7T�+��O}",�ʵz�q(�ks�ԓ��.\\�J���R=�qL�b^V1��䓊j'���+���CjF�+F��A���\����k�u�_gJ��7���j�R���k�^��ϸ��:�� /�gU*��Y=aw�[�ԬY�r��IŦѣ�7nmnj�i�O���2�4f�֭[�X���^{Zr�?���y�����5[�ٗZ[!���&�l[��F����-[p*�B��̢E��^v5��s�e��H��[���y�{��ɭu�������o��9ں�W������o��u�m}����;�\�C� �_nn��8�i	Ç�ظq�.s�d��`����3f�0� �RZ/��2 ��1�&���Иҥ� �P�xi>���m۶|p����׭q�{�zU�����~����P�������^��6����w��Z��}�����u���D^K� }]!��GW��aÆ�5�$�����A�`}�w��ׯ?�C�X ��nݺ�̙3g@�΂�H�&t��g�-naڳ�O�3��9�Qc}�� �?B�j>���7����^��|����V��`�������)_�J��N����{������A��ެY=� ��� ���-�~��A�zR=ަ$��y�����rl��QO~�{��5E����wUX�:C�~�?�~��+��+}�l)��$� f�n�*���6��ȣǏ�g�:@�׺Z��t�k֛����t0`�i�g��:Q+ʉ㇏�5,�ܼd�#?�z�=���>������4�:z~뎝���+G&j��---C��.�F��Ţ7R�ut��HxQܘv��\���iU,<UL�e�:C�Έ\oF_�?Sk������SEk_��W���u����?Uy5�N�R G1pd�җ�{��TJ�M��5u�T����I^z�,| �X�xqkkk��]�7v��8I&M��~����$Nڶ��r=qɃ�Ь7*����uQlekݺy�ގ���:�3q� �nl�^�t�y@������Q������)G}�����1���>c�����g�~f���2�3]�`��	���ӑ�?��̒�j��&�3�s`KXrN���( �������&T�ODQ@��AI"6�,��8��ir����o�{�Psg��]u��}����w�VW�:�=�N��S곙ơ��Ip�W�\`�ڵ�r0hРY3f����*�V�Yݝ�=c�^����1���Is���q���M[L��P����vP��!n����S�����#z^�O����쓨]}��<�3᧑���l�t�3,zSY�~�3측;���yS��歫��'���0�:{��>Rю����Ů�v��B�h;8�c�L	~���w���B�]���uuuЌ���#F���Ｔv�+�$j����5�U&�}�g�MM�>IV]�!��{����c����'����_^д|yvŊ����1�o��$㱌�ww��֭�ܠ�H�y��(2����/�3�^�gy��������?��;���޼¿x�j>�;�]8���,����6a�32���5kO��~yy9O5@.<������q�pL������qy{��lN���Ν;��"d�GwU�t�4�k��X,H'�z�B�������}�����a/�?�g�����q��A^���L}p��P__X?h���N�L��X�Tb���U���<�Lg{��5k ����lٲ���d"�Ҽv�Bs����i'�ή㞾���x>�\y}sJK_�������rHQG��n��mj���h�Mo�*is�$U6[5�9�b�7,��2B��]o�����lԑJW�Y/���w\�z1����z���n�0����1�NBVQ��$��2ɸ&EAN�ǘ�Tfa�������<x�����|Pb˖-�t���V�;ߤSw��\S3�r�.^u�*r�͛6�שtSo��V�j�<��7��բ�0J�&�G�EEe�L.���L3�8��f1=�U�\���W>��.;K����n�k� �g��_���?�o� 
�>�<�'�I$��FaVC� �)O&����J5>a�d?k�h_�t)��֖�C���� :�؇z ~��U� _�(=f܄����y(O��3�����y@E3gΌ'RA�$�R72G�<{�Q���ϵk�]mc~��*�ɤc&�p���7��+++w�1}���S�W��Ҽm���e1�O7����a��iSw[���ŋ�;^���cF-ysK7:Y��x���������3x��Lw�ZG[d;N�f����hS�Џ̦���{]���t��\��x��R?����Q%�X��5�Ϛu]5]R�e���l��GA�n��STtK�_Ɂ������-}��Ci�S�E�.�5>=��X`����t-�E��O��f��U�Vis�&Y1u��a{ͨ������y睹/�XYS�li���������ЕR&N��p��|��I�w��q�V�X�����D��#f�G�HJ]��4T4��|��X*_�X��/�v�����������g��
���T��ս�`�	��d�2H�n��ƃn�#˗/t������Gl����+W�?>�Gp M˗��d5�//+����ꃼ��U�HJ�7�G��ɟ�۹p�.J�|Ϯ����u׿�2��}|�ꫯΞ1���m������]��UUU�G��زm�o�ٶY�v�k�����Dl���KV�����w!M�X�رc��5�O$�)�A�֭����q�0�9�O���J=��������	�H(�?�����'r�nm�'�~A���t+��t����M��͍��Q��KL�w��ʶ�D�"����#]��e��DP#Ef��<.�v$�a�qX�bS�|�?��Y����;e�4ХDtz���*�*+Y�/�ͬY�4����e�^����$F��v��͙�^��L���v���e]���mЕ#GN�c�X����QY�_�n��7����=�Æ�:�����ڙaŊ��[���[Ƭ����ˇ�L��Qm�-�{"/����l��R��J� f΋Q���y����s�a^ڏ��$��Ev�����bW�;�^�Os5 ��푂Х�G��c���,Bi>������!�Gy�%��N{�X�N2�!ӛ]�f-�˄	Ǝ	���ݩ�`��w6nܸb�Ҙﵶw�^�a�!Ю�&�߲���M�Y��v�a��Ty��'�9z�^h��e�ΧKF�t� /b���)M�]�ٮ��׮c�bW�~�z��Vة���!���+�.]�rՈ#F�L��s�e����28�,A������5q�1c�ԛ
乌����iÚ5k�h�hѢ!C�4ԖWU����ܬ�e�^<��;]t2f�t鞂\M3]E6�0���h�%�v�>�"��o�]Tp�����L@��~�.�|��/�AK�O�Ea�o�g��l�
��J����V]�Qm��G�nk�W�M5�BE�\
u����K�'�[�̽v6�Xm��UL�v����G�-��sɔj2�%���3f� p�j�A��������@*չ�!ӱ��b���Um�lGG�S"��ٳg�*uT�Je�#����V�T��uū�_٭�2&M��֢�=�ܼW^�R�(�v����h�1����
c�kU�qK]{4�ӣ|��R�y��F��#����1������mg��W�?���㮻���r�ǵ���s9H��"��	cu��-k�tz���ʜ����C�N�������?���1�ȸQ��nc�i�J��Sٞt.K�"'��V^� �$�L�[�6�8hb�����d���������R�v���b������\�'K��\�'�>��C�@W	� @��-c�0��AUC�Ĕ)��p��իWw���3i����--��Q<�m���w��r����N/��eL�Uka<[p�d.h��Y���a�Y=�^��p�O
~��1wѵ��|g��~W�i����T����_1�+�ٔ����b������T�F5ʈ�9�ׇA<Ud�]Y*�'�k�xJW��eB݁Ҥ�+?iZc���	�~���G�f�-[��Z�jݺul�5`� ���I�A�/tdJ޲�<7n>ikk��}�7XVO�=i�����;��3�N
���	08�5k�2g�?��	Ɗ59�w�.?��&M�8r��d��ڱ�yɒ%�[�nj�ԙ�)4&�G�#UV��Lg�X,�➊'+�w'Tֽ��k^K.�ۺ������U����e���ľ���g�q��a�C��l�45V�7��X�,��E�#F�V��Nj���ޱ��|]�PuᑃԠJ�'���t�7d���*�[=�a�СCfL q�� ��ܴiӒT}l��Ԟ}eAӺu	�:z��3=��~��t�NL1S�H�U��d쮅1�L���dgP,L�ʕ+����:��]Y-M!�ˏ���,�������N�>��.Лo��q�Fp'*��B��+~n����Ւ���<�K@���������n�+�n��ـ-��l�߷��4�K	��5�L�4|�pvΒ� sJ�9��N!r����$��'���18��s� �n����A�m�X�K����e36���C� �z{*1a�?�ߺu+g"ė���=dON���d�K�O;k�,�%�a�6,\�0��7�ѹ��3�ga��WU�f��X˖�k׮�1�=�r���**�_�\�<gȐ��C��p�;][�۷��#TaX[YYk�Nb!6�n��7�o������Vk�Ѵ�)����_�q�(��,�>f�%M�֠?Ooۚ5qJ��<�M�`O����O��ϓ��Z� �& �������@m�.�����O�J��>;������DAY����'OC�w2Vzj:��m��I9���ma��Q)�Mf CB��M��������1�����.���*%Ĥ~9߈���3:�4ǜgϞ����v==�p;��,L��hJT�f��"�ga}��Ǝ� ����oc!(q�ܕ��r	H��v,�0v�c(��Y4�m������u�A������I6��l1m0<~�=
\_�����E�Ü%ӽ���'t1�0�ܹs�@�G��AO�<���~0�^�E�|2z̸�k�U�W��uN_�7�0r�V}�<wŦM��~���C��9`kk+��w�u�Q S����Oǻ�U��aC�����l:^VX�7M�L˹0���3�$�I�o�q�E���194��O�3
O�Ù�yO�*P��%��4�*s�ɐ+���r��o+Yl|ezo���-��dȢ[/^�
��v
�����*]M�g8I|e��G��u7�T
4�C�`!�-��pG�͢t&f�k��i|+Ɣ"��܌�������p��)�{g+����"s�4��!S�)XR�&�y�B�uZ��UA[b�'s�8q"ǴA
��i�i��&؋�.XMA8���@	�'�F�b~��t�R<(0�Q���̱�aH�V����wm��}����.��`d?���^!�4<(c���PX9葏}�c�Ї`�u��JP�`�,Xp�M7͛7��;H3 7V*����y��m������z( #���P
�ׯ�W~��_�)��/h�V@b�wRY:�^x����G�/��
0P�=��o�[�>g?�zV9퐸*S�N�ԧ>5g�@�	�٨��а/<��w��������œ^.���ӛ������
�\eE�^��oեCh�7�^���bŌ��j��?~�ډ'�pB�!3�j�����b�l��H�����=Ue�Y���@��v�+���>���舃�;4��ui�M5�\��|᠃��.����=T-O��&�̅��v�m�o�	�wuvJ��o:"�*	�I
9��'>�я~�|��%"gO���'���ʻ֝©l�BQӞ�VÞ����|�#�~8��c�@��_�~饗�j�h�"ͼ(�b��!��җ���xx�S���o�������D���a�2􅤝$8m�}����?�����HP[�|ٲe�u���z�"}y�]/��D��gQ�|�<�S �Yי1k���Ux���z�ږ[o�}�8�ƅ���$|���������?��;�����f�"�P���sz���`,��`pxt�-�y9�x뭷~��{�9�c��gθܺ�N�����r�!xbgC#�4n��^\h犊O<���O��֛bY$8h��-Z��uσ�FX�lZ�|��`�ln�L������:�N;��{W����/���`�L����[ S���yl��l�d��Γ?ic.�	Ky�9�ཆi���xA�L��OFN�4���z���|Ɋ��;�<�1��W�
�����O=��Xp�r:I���J��_�.����>��� �fƣ��<����W�w�qL	Bn��S��1�I'�UC!�I7�sP����I�y��tHl/jY\ řg�	m�O����PbPe�6���Ff�<�
�=�e��s���^P��c�6��?a0I��^x�[n�&�U�P���O$<�(�<���S�PD�߂,O?�440���V�v��t:?�����c>o���2[[�ݝ�����;�#Ə��UW�*��a���ګo`����Eh>�Ep��5�	O锂ߠ�@�:C�W ��� ����+�K	��ںKF�
����`��������r�Ygv�a�A	X /� �s\P+z�+�g#ap�9 nǻS�b)a��.~��@Ur��N��J7T�2�v�駃'��x)�U1s)�n�c`=%�G=e|W�$F�n� ���9s&fE'��z+��Oz���َ0�}�9&�\���3E�cp��� �7@	�s�;D����r��f�ݶe"��\*O��b��EI%� ��@�%n.���_�,VF�Q}A� J�'�f͂������  ��w�Ͷ�`Ti���i����	F%�'��W��w�����7�gT�td�ӯ�1�̓0�>�W�)�T����bYOyA�5u�(�p�s�a�Q���'���j.��>��c`�A��G_7 ������~���������N��ӭSB�\W������/|�.`<�o2a�e���{>����.�_�/N�I��DX��V����>����d&5悧x��+��̪|%�3�E������KAL�OcX?Sᕩ$vrȨ���_�|������k�]�xY<��d,�����ѥr]�����a����YL~���i���� O��
t�viN��f�*kc~kN͘���a�e3�<x�}��6�V��IU�]���b�%Z��'{ؤ����4`�[;Z����m����v���|�r����*��C�&+��� jR:q��}���q�7�����;�1�3��u��lN�aP�£����1y�	F��r(k�&���!�?���ˑ��i�Mj�D4~��;�䓿�����Q�J3�&�L��S�<�^l%���y�:�l�K.��;�A�
 �w�qNp;D����`_	��q�	9����W]�� t������}�{0?P����)�^96�(�,���+���@�rӀ�H�l���~����]vQ$	���m�������F��i���s���+�E�s}6�ׁ;/��bL�j&��f�����?��W���V��B�V��wv�%�]���2�܀�"xB
K�Ebf!���O�2�t�MA�C��f$��O���1�\�F �����p+$�{�9��x��w��7�[���#�_�Zn(�SG	�����b0�ׁ�;���o��f��͛7+�m�P�\�D0�x�8����������n zsa���S�Pr^�K��\D ���ӯ��:��9z��9z���@|(�?��(V#C�@��� /\_�`�B�~!F�bp�#X�z#pc
��%���=�я~`��5FF(�^������X�c�=4�馛\��r�c�(.8��fC�c:â�U 0ػSO=��_�:�FV�b��)��ӭ���a==����ںA]]�H�1������J!)����
<�O�6Z��{������F���րӠ����e#*(��_��W�0>�ȕ�" �� �����z�,P^��U�U\f.,t�ԩSK"Or�l���n��0d�.��׷-�Y`��s��"R|x��� �@I���?���wd����"�$(v�W�r�)�"�g�18�l�i?�裔#jH�����W�W���78[ʈ2,��a2����_ ��<�ؾ?��=s�\�����Y)O���+ܼ=���l��r�$�k*��}��Ӌ�w/��c�9�/��4Hp|�p�	'|�߄k�R=󢽓�M(����j�}���+���S wX���:�g?���l��FZ�O�����������v�&o�C̅�������&�wU�� R�o�4��	�������?�z�8���b��/^U�7�(^�L?a��X`Z��YʻI:���<������!�����F�����S �<`!�,�-���kb���^N�]?��B�ʘ�SO=E�=�\���8&�/~�3������d2?f <��d~2J������^���7ޘ*dH��%�]�(��R�� 7��k׮fvigt�58U�gutv�s�o���#�UW�� �u�І����3�4rg���V��#M�u� U������زZ���=&ȅ����T2PAyy*�I�9mH�9��A�:U:�'�5H1�M�ݨ3~?��a����D[Ȩ�)���'�y1��^{��K�P��Q*G��g?�Y���E���e��"�aA@()��DT��8��%\�12��h��̀%�X����a
0����0������͉�i'p���p� @u۶m+�����	�	90@���'�#���m���V ����ǅ�3����\��r� �0��=�6�`�ʕ�x)F�������`��&���/Dc�e�n��2��������B|��5����N;�����x�m�(�cQ�۫u=T0�^����3j$
#�SȺ;1�q��� t�wp��7������O~�����NWF�sE�a����T��^�KIJ!�]�l���_0���1��}��[�lA:�ƻ��)&**��Lj�z��w����۰�s]���/�?_�򗡠�6l`j�3�wc�����f�	 i���G���*���%��/~�!WHxL�$�(�߂ng��BU���N�'�2H��B�ͷ�g���ٞ*1�2�
�˸,�@=On�m ;pV
w���[�p#��#�y�7���j@@�x�y�b��1c���'@jsss�:z����sL��f	���-�� �����2.���͂X��[�x����'�fM/����x1���X�]��g�: @Am��'�|������ .�"�/��2�2�a�&�/�=s������K	j@ق��r='Q�ds�q��O?<�$=���iM@O�#�)���"y�$UfW�?묳(�Pֈ���AhiP 2K Aq.���"�
N ^�eZ*+ɴ���5������XYJ�]�畵G��2ۭ'�t���L+�1u?� ����_T(�6�V9)Yj �����$14o �S$1,n�Or;7O
&,YUD���Q�6ԋx�܅����~�5�\�������.�d.`b� �L}���H��>�[h �t��y��q��r|�	L��@����r3>��'��!M@���S;߉�RJT�FxY����Fd4h��Xz��D�fc^)��<VV���k	�[��8�� 9���եLR�����.�S��<��+	3`<�i��ט���m�Q�&j���TXnX��D"�䵹�z�S{6��Yq��e3f� ۝|���V�r�y1�|��GC�Cl��`+��+%���Ga
ZIyڃ�H�I-=� .�����d�l�$R*�n�ܺ�99i�Z�������1|�����<yȸ.�1͔xU�_�����U,�����ڸuKWuM2���EoY���E�w�}�Luy�1��i=US�j��.�e��T�^���������C���T.&)h�T:P���FB(��.�j~�gtr';V�~Fy�LbD�r�W vKH����R�����I�6�F�Evi`�'0�  �y��N��*��$�ݘ��%O<蠃 �T�0ZL��xj+J>f� 4�g�O4���9�w���������>���I��j����D����e$�$�a�~��9s�PcRܨ+	������ch�U�V������aث���[𜭲�Զd>�� ��
�)Ay�]|��/�Mc�Tl� Ɖخ��{Ƞ�/�|SӺn�Q[�0P���:`�����V,�<u
>���P� ��\�?���L'���1�N_�h��ѕ?�ش~��C�@&܃�&����ʬ�G}$�H�Q���AAɀ"�����g��'�[�������
Y�恁���c�`xKZ8.1�<�s���8����ᘘ-��.��uC$d0�U2�O��nڴ�`3ǳ9K��	f�T���s)�B+��=��Up�7RĘA��hq�Q1T��re�~Ѯ���\	�����k�tEN���N��~8�g������&�y�;�5T m� Q�k����O}
d�����$�����q�޺u+D�����:;�"�1h$��c}Ĥ�É'�a0g�vZ�|���[ZZ׬Y3y�dp����׿9hP^<���e��;��&"k&M���o^�|�R(a�0�^���x<|a���K�,���49�A����.�L,+@9H$@&�,��?ْ��p?����c�g�]���%d��_N;�4�v /����\�����A�)�q� SgҨ��/~�X5�N�$�@��^{��,
��C،+ˈ�^{�ݎ�{�W�q�~��d�q���ǎK>�#�d�z��.�Ja�\p�6�Fsa�{��``�b��Cf��De�)A����l<�� ��,tC.Ll�y3�Ô9e5Ld�a�9���}�k��c�=&�(1~�e���s�=���jh RU�T�7��F\(:�!c٨����)�rI|���x�3�8�&R� ��ݨd���Q߀�����K�����<��yA��L�9P
�t�O�-���"�!>�?���o�]YI�`�?9p3HơHz�M�	���|����<2 ��20l	p�H���r'a
�/��N��A�����6�ϟ.2�5��(tn�(��T�ޠ��m��M"�r����@p���1��:z���3��Y�~��3)��Y�:%X�e7н�BU�W��m&�)][�ɜ�A���# �ǎ��km���h���M��!��:�{l����=�	�������������\<�Bap(����G&�'N�����m���H(����%�L���?���ĺ���9<b���Ъ�w0��<88�3X`S��~���￿X��U+��9s&x@�64!��";�c����^��[�6
O����"D�@�t�.��b$�?���+,`�_@�r!1*|�%� �3�,�&�E)p��a�)0y�(M|������y$�D�*wR}ˬ�����z��̀����]ĝ���<�h@	&`|���_��#�v���%�`xp>����%�2ݛ�wwuI�������ú\z��C�x�	8������qyH����֭��S�����09�(YT9�Df�r�}��v z�ٽu��Κ5�N�p]zb.�0܋�b�.\����-9?<����/"��j
\qS� )���?��Cq6(��@	�v���W�3.�=�������3�.q�Q�9ǝ �9{��~5��S�:��ռ�˰��q�Y]�?�?& </���-���N=��7�x�$֊61pNA��e~�x;H��FFv�	�u�Y���^}��brDe��Nx��)9�T?G���4|����W��j���� ��R+V��0a���a8x�������toF��d��$|����������[ZZ �u�Ux)���/]�tժU�&Г!EB��"�L*�w�M�����ni��s���4H�����Fh�&�{���̓ngj����}��<��>���&��a��bKF-�� ;�H��g�.�9r�(y�\��ԩS�഍7���r,y�_���{3G���������QG�W��?TV��qv�Ǉ�a��Yy��G6��Y^`�Ȟ:���O?���'����l�ɂ�
�C8��̷����.�<��/��(O9�_Y�!���Z��+W	(�����o7�V	�TB���-�����!������I*3���O%�a�*���^�Ky��tYϲ@��d�Rk���Td5��#/������)5�grb��@5̙�W:���&gH*�E�������!����_���1�udc�	te���@�<�@��+�P�r�
x�
�ՏK.�P��z�p������)�B΍fe��`��x.�U�|� ՙ��(z\��"VVQYqΙ���[�mU5��:�'SYQOG��6�vά�\����F̜0|X��oS,�H���R�����X�Փ��Vڷj�D��WmΫ<�39����}[W�^����ФB=�X͔�ds3���O���m�J�T��r*���L�I&|�O ��Q�{>hr�!�����T���<��Y�O<�OBY�f5x�V��ZD�y�i��w�}P��8�3O����]1�"��ߓU���/���Bq���+W�P�$�?�&N���JI��PQ1t�8�3��]w�%Ņ�!pJaD6	̒m.j(��ge�#��6��=W����R�O���d�F6'R$��x�I�i�N�
��x@���9��G�t�I�v��)�X\:�M*��P� � ��\/��O>��G�2	�p���.�֨Q�>���ޘ7� ����to��H6��?��U5�P\�&M��C8Zo��d'�<e*}]
\g���߅zF���x�՗��cF�tuu0�H��.ܕ}�ه6�w�i�U"-\`kk@+B���Gvc� ڒ[��X���2�(��M�6�,���y��z�j�����Ӄ�̞=;t6�5������<�.�ݕ)��ȑ#1��C�*��so��Ji�"�w�����G�܂P��`�)��"H!���p�-�q�w�GB�Ha"7��o��A|x�����e�h���+�=�/��;�n�`���Q6 f�P��9u�*�X�I>�,m�1�h^R�����}]!����ٱ�{�7��%#&l ���qC�V]�i����B�q����4�~.��(8,���{uu5==i��}�ٷ�z�>�읦� ��hm	�c�^�-dlj]w�}�/�_��/�����땓8�EӃ�9�裡���L[�##�!j?X�{u��)� �Lc^�$��ZȞ�R��~0_��W��g���9�Ɏ�����Q��DXVZme��Dɸ�Ϗ9�7���3�r�!s���\�$�C �x2�Y6�/�6�id�s)M�|��o���	�6W�]D��`@� �FG���K榉����M^�<y2��/~�ȹdp����|�<�:[���%�������o����~�r�0�3�v^k�Q�x:�. ��+\����W��h�5���tڨٻ�Y{<��kQ���t�A�,��ݍ`:.@�;�*�w,!�h�"��vߊt���i.����xnЂ��;�S �I#	�t޼S8``@��8�����ypp�| �x
�v`T�y��lNr�p� �3AW=��C]�9��= _�%Xk����9�/�k���b��twtu���:��fBxyU�X��(Ĳqp�ٍ7ވ���άmkkj*�����X�Dj����i>k�(+��ɪl���4j�ipO���%{�(�x���C��ӽ�w��rVR� ����g��[=S�����gɒ%<���a��q����%�Q��-u���׻�/�E$l���o- �~8�m�8�
���od�<�|��g�Ⱦ�0<�7s�L�E�F������'���N�'����o�ʱ�g�Ϡ��9'Fkd��^ܩ>F�(�'��Q�544`��cPҞ�[._�x&{��'W�/��0���T��u��k��Bü��k@^*�'L�2c���'�`], �-��y�
jA�$0u���#���Ig�5�0��o�M�>�f����y#�7�j����bwe����J?�� � t��X��ncc#�h�C7��u�
Ċ7@�B5mܸ�9�(���p��yYY_�K���dFA!Y�<�����ۃ{�$ɜnd��QF�s�G8�z�F��)��ɚ�2C��v\����Y�:����E�(1 ��澊gj�0�s6+���{��p#ޗ�C\be�g~n�{ｙ%���F7I�R�I�F�/��R����/ē�����ʦ���ꊺ���>���>}h�@em-���Q�֭[�ʖ��L��D�aH@� fIw����a�R��"�-���o�qЈ����UvA^h	�d<˛3��]	[��y<�+9a��N�f)f���0�t9�r�(�+-���5k�s�=�Cëu�Q�����_N�r�EQ'|�#�馛���t�E���#��E	ҋ �=�J=�����#��|_Xm�D6=r�@���+eŇ M�2�g ��`<n![�y���ry��sʾ�	|�(j�k��0�l,�st�tܸq�J�������tf��)D���m��p���I�
�|_Q2�*H,�{���3�<����v�����VS�~�s�H0���"^�IP�n���gb�՛�u�'��d�������u���H+��m�f����>��_X�+�z1�� 6�T괠h̸�&MLhX�� �-nm�Q7��A�_7E��~q���z��w;��K�^\��=)M}Z �埸�P�fS
Bey�2g�����mD �3m�4wǊb\���,�24���c�_&�R������O����c�O�����[S��j�֮ގl�a�h E����N%W��0�)�K��s�>O�PZ[�ꌩ����W������S?������Y�����
?���F�W��8poU_��I�JeC�LJ�+�J� я3U���{Έa×�wY{�'��%B��u�O�=~&2p}E�1q��Q��U�hcǎ��bɎp�ȣ�O�(��o����䚒+\��������#琜�)���_x,֋/�(����T�|)�s�c�XB^n�R�X)���r0+p��Yt#L�j0N<��Ҽ���8�^0l�G�7o��N�8h4���S Y�@)��Psw�yg1���;pN�o�Ũo�Y>������|!&��ohЬb��/<aJ⒥� ��60(�Qu�O;��rё�fzM�\��}������cta3�|�.��0t��I�-�`���t�B�!
���a{�R��� �^Gp-����p�^��.:h����
H
n~�A������6�v`�����C�ܳ�Y�������r�N�D[�u����	�>eʔe˖)G`����'�2
�_��3W~AL v���E ž�ΡC���*k��}�I��"&�/�s���+���*[�Lw�;������WF�� 8��_V}C�B<��u2��\Vt=4���:܌����v�Z�#9b�nS��vuCb0BGGGg{G��V����G��3"�i�ꉪ�#��c����m�zᰋ'V�8�\.3�t?>Z�Mͧ�~:׷?L��󁞁��}��~�J0:��B�^x��!�t�F^j�e�l�Fej���AV�������i�i�����ܤ��'��|X �hr����� _唟w'/:�߅�8��o��6e�:(Ǘ�m��?n�O��
�R�7��0g�8sN���>��������$"�%��7E{�a.\��}-\=�gA�&�y�h��Z�n�0 .� cƌ�_-��)x��0w3�������DH��X�T����k@0��N#�nէ���L�֍�6ll���[�:��$|��Z��s!���s�K@�j������C�y�ȝ.+K�-��e�����4R���S�.$.8?Q����@�bnܔ�?e�Y��6�!�(b;?10�>Fa����l����2ٖ��L��6��}S�}��Cy�/T�\�D���ΞN�v:��~s�I�4'�R><�|Y7]4��B��[A&���-���u�Ad}����ЛPRR�Q��B�&��&�r�K���x��`Z��c� a>#y>%�R�aS���k���^�Q�}`�S���!<#a�]#<�$�&l�p�e��v 4���	g��y}�^�%Kc�G@NC�=\�*��d3��C�e��l���p��]���_��0+p����Ap`���w-�k�ĊP��<<��枼?�����d�mۆշ16`}�:>uLr��(����gxktΖ�	\}P���ܕ�OX��Y�Zs���*�̀���qxzܖfR;vy�`�D�%W�[�R��F`´%�C�`3߷�����v}dXw%�XY0� $	�1*���e���^<���{m����1��EPl����S��"�eQZ��f�V�:�����W
�*���n��N���)8U����|�}/L���Y���i�	�V��5��0y�V��LA�r���J���7ٿ/9��@]GH�p�$�I���%+��:wcJ�.re	QXB��>�l����X��g�s�-I���r�.f_�k*a�P3w3 $xT�J��08T�((n�7�3����mG������P�Tܒ�Qd�@w�����]�㈡���L1ax��r�O�~�Rl��_��efX�Z9YO��wŠad��Jؘ�0[�|iȐ���bt㾜g�^l���p�&Y�����Gmho�4$UW���T�ccj�Vaɭ�
l�eu��D՚��ʺ����� �`CϜ	��8��������r�"���&3@2Ŝ�/�TjV%K��^�S,�Q��_�t�r��9�5���rs	gȴ���}���:WEq�7b��蟾�e<�[���z���AA*�zzcal]��1z���-����/��T�~�^�f��L'ksPx��g��J<"�i�S/�%�{6D�b��T<橪@�*��L�7�#8٘�^�NiL%��Z�,���\���K��XD�e�滃�K�G!T��憗o�����G<�XpQ��y��Uy(��N�Adȼ�ݕ�EP������DR��ԥ��k2&�F)�9���L�H�&��P��'�S%��r���cU��H6�N`���|[>�����^��.8�Wp?=�WQ��xB��0D ��-eɔio�J!2i/*�Rۢ���s�4���Kx�$��qҽ��IQ6F^S|x~�*K��A�{Бk���������Й�Z:�kſ�������3	c�k��t�������_s��хNǺ�9�����2�����5��M���b����w�������0Ӂ�;�/��K��DD"�Ͻ8��_�Q�8��P�yV6M(���;���`ڒ�*�Ul�2��$a�Y��u��|�9����VV�y*�#/��8�|��iؠ�r��Rř�!�.,\�ش�x�&�.�V�ZL�/T(v����	;{��T���%���^i���ĞJ�
s �U%�Tl>^ߘ:�MR��L0��)7���:�%���� ��Ȟ�U&�!��I�.1N �e|h`��s�|/23,S���J�&f��o�G�6��ݜ$��%�h"�|U߬����LNc'5����|r���������� ��t�r���I��FO�&��Δ�,ׇ�L  ��IDAT�P~�)ۢtZBce#Z�ŘZ���;z��):^:�/�g��eE��&��C�*�"��,R 0�zdE&��s9��a��]�#J���%�����Xc	�ry���x+K��@��J�B���E�bgk{�� �e>��ű��-[���XvP�$M��ػ؂���J�*U2���>	|ݼ���ڸ�Z��
�lJ�(��G+�ygd�~���VT	�D��:����BX�lmm%����^�SђP8t����
,4~vvv��XB�u��v��m�[01���0�w)�@hBq�5*),j^z�EY�!Y����ᶂ���v�.�T���e��FݘN-�#�ʞIc�k&m���Ç��ձ�<���)�	�e˖q5m�/����&�cMR�Ŕ��
t����>�eq��(�pEi&j�&�`e�Ȟ��W]��
\#�S�Υg2J6�K�bOd894��YR� �o�G�|(O)��2��x�l-*���,��잌��T�"ڌ��w;��%�H���tg%B��[�n�g`��T%�%
�R��G�^$o�)��S
nBHs�Z����̙������,5Fί��i�h�r����?_y�>3c��)��`�m|�����KT̩~�5�b�6���Ң�?ዒ"��Y���[����#$�������S�y�%�/��� e[��c��/��]׈W`�0-��8��� �N��,Ai�����I=)ʙ3����Vq?��8z����E3ʦ�d�h�s��Ĕ��}��\��;�|�6 �M�U�JP x�`Ǧ4���š�����)#�ӓNh���$�M�)�'�+|�\�+�k25�k�*�6��kD�q�C�������k����0��xѨy��Y�N��E�%�[�]��������iOdh��b�jiiqo(�v�?���q�F�h�o�4W�cp,!����>f՝�Y5���NR�U�6?�e֪Ly�|],[9}7�a:�	��嵙D&QW5h�8��޵�y�?v�n�9�]�%b=�j�M]E6�J&��1?V����kx��5{A�'�YӴ^�yٜ�vJ����?#���D�oZ�1ە��4'�%�4ctЊ8�X�U�V555���5?w�߀b6l�	)Aj���+�y֡H�4 �ʕ+I�������ߗ.]���j�@�o�477ӂ
vh�k޼y.��bR/ݼ+V��Fp�k�@�d�����wP�ċ��Y�D�*�xe�]��%,�eڶm�a���Q�f�(��3V$�k���]�x���O�L����ωǓ�Y9���Y�����SaY*��-LS�)�˧<d߼������=��w2�T�c�66K%�ɳ�V�ǌ���a^�^�w���Ǣ�����}� �u���
'�Β%Kb6�~�T��T��t�b�xh�3&��&Мwb�xB�����%\S���Ieqd{3��[�nǷ]��e�^�g�L�m�4���=J_�S���ENgS�ɲ�AL��R�q��;h,��{)�������ak����r1�t	���[[[�́�kݲ9Ȥ��� g��U����޺m̘Q��5Tc���ԞF�W��LL��d}q]`�[[���o�Ҁhگ��垌gs&K���OnT%��d >H�J�G�A�?������;�m����"�y��ׯw��0V7xNu��]�s����
�i`'#��Hlp+�ێ�k�W�c��}{&���uA�S� �Ek62d	�WN�-� K�aR"�+�~[)�q��#{0 Y&N�(�� �aL��ր!i��իW� n���t�h��Op{���x�2����*mN�i��5���9Υ����G��B"�Q>�b�	BhHW7(*�#.���������.��]��{p���<|��\�{&�z�Q�f܆aa�qdӹ����d`������'MƎ˕��5�0q�,�v����(R"��R�^xgN�f!�ӧO�f��ϲl�Z+��հj��)�:��S鱄�ubMyYE
�@￤L���0���ds[�]��Q��tj��a:��3��\��P|�7�xs�g�(������S �#Ν;WΧ�g�Rb��t0m�/(^p�m�<��񳠭�{���9Ӂab�꫏J<�;��_i�
b	��BC.���eK�H9���T�@�䟁i��p��c�=� ��x�j-��y�1{��}&�CܦL����3p��a;��c�=�-ުZ�x1��J��u]`fԐ� de%\�4�	,1�3g��=�wڰ�^{�M��u�kɤ�#G�+Ԋ�}��z�,��&�=���ە��^��_��xe0�Ur3~Yg.FT���3'��.!/  4ưa�"[�+�q$��������Ί��ꫯ�L�Z�^�Ue�
�:Ʉ���x�	?xM�	��ʂ����4d�6m�v���­<���'�t��*��72b� N�#�vtv.]����<�L��g���7�?�0�;\�&�s�0bd�w�OoΛ��V�o��1� q�g��4@������8�?�M����fS���o���],�	����C[�D���ב8���_0�]~�n_�7N��z�:�q�s�=W@��W���T[zWA��S�]Ͽ�9�Q`V�*@���#��s����1O豕+W��1�R����LT�N�.�:r� �6�J�Y�����*qp�_B���za)���e�Át�Eww��~�Ĝ�d��z�����1�@�����f͚��O�9gN@:M��+^Q�����D��vVT�������798�a"�����X<���R>y��y�)S�C>���&NM$��5C9p��/��Wα�w'jw� �@fGydh����O)��Vx��G!0�n�<��'�p3��=��9V���wZ�/�Gy���Z����t�[	G7ʔaL�&�� ��*Y���ꋶ6��>NZ<���[���kݦ��T��D*�|�Jp�>���zǇ�#����D*�ˆVfC�Pd2�c��)�Qy�O=�~�J�чz�Pܨ��>�v����z���X>e�T�
���+S2�h��6H��Ĝ���u�Q;0�lb�1{衇r�z�; 8�p�)�R�dRP��1��K��I��ПQ<��Z��*i�qP&tdP(�����H�!�R��h�N������OM�3�i������SOd)Av1��Iss�?���c��y��0�X��;����Ί��s�Yŋ7��=X}�L��G%Z&kټ��-Yn�]iܼf��捛=S�n�^{^@�EAXY^�Q��b�׬Y�St��5]]�I�,<�5	\���Zx_XzҤO0rʴ�k�h�a�����v��2��8����$��M&N��6",}�V 8[{��J�Af��ٳg36/S*�)[	��7���Jت�	������}����.�1�������"��������𠠁��\�A�8TY�?�Wb�+V�?����C��u�6ןk��*�D�d�o�) #���� 0�n���W�߳%�^x����{����k��	��A�,[s �x��ǏUA�g�u�r2ѥ��֖�y�]���X^��!��m���
#��7�|�Q89���dM#�T*L���PV����y��0k���9&����zjΜ9�M-V��N@0si?��H$�ݮ_�,�{AL�9Q0y�,�3�/���͂02���]�e�p�uuu1[9Z�*����lg1���c��>�X`��#�B����{O`���'�qi�݋b?
�$(q2#g3�����c�:thi�0�u���}a�K�g���v��I�&q_N��Be���3�dF�iʐ���Y#s�9�Ϡ�(��p �]qGg����X�aG{��?|�N�0q|	*N�
�qx�<E�fnJe`����;��{o߮G���?���~.���/��"���Q���̈���3τ�[��މ���r�)��;_w�m��b�,3!���[�L��ʯ�):/k�A�2y�[o��g���*��Ă�gΜY���^���J-���]<{�@�x�y�j(�--�b	? ��T2�29�a�OH��-X>@[B�A*�@(7��a+e�u���y�����s.D�|^z�%F���,7
���m0����%�-e��`J0<��X�"�M�3Ψ���)�a�>������$l@������k5��}��?=۩Q�M��h/X���7ޘ:ujT�^���Q����a���Y��=�u��=餓�㶥K1:p	���GYb�@4(��;�E��a(�ɷIM���������TS�&H7$����v�G���s��ǀi �^z�ه�� ��e���H���6�{9C|��d2X�s>y6- �Ձ^0<pa{��G�|$]_�/4&�2�j�.r�m���F��n��O[[t�9���ឰ*E�����!�����	$^���[o2d��3ٮ4��e���H��hp* �v��C�K2�DC=g�
k����?T!��?mٱ$F��J�[��EV��D����= "�X�yƜB�X�6��̜vѿ�	������X:����t\�~��1, XN3y�n���<�|[Q��O��)�$g*�WUUf����>�)���l���[@罽�q�����r@�x≓'O��z%s͕��w�y's�ܨp	��۱F@�#F��n���C���O��y�ܾz�jH4dCC�lp{�a��[O5�=w��=��S��L�ؔ@��˗3���(��Y�p��N�>��]
���	���{��?�x)�6�9i`���-D�ʐHZl���|��^{��A���(AF�@���
�$�)���+f��<�����f��j��i��6|�pIH)62�M��v�����&�W։��x&֣�2z�n[\�}艪��������k׿��i��N
�lN��x~�w"?й=�����?������wU�3�����Y?�i�h�$>�'�+������
����M��s������%�EE �t�uׁ�Y^O84��<��;����8K���\}���֥t�{�5'���:�1ˌO��e+����?|���oh���T+�:�*�ƓU��^�n\�����ƺ�i��xqE��+�[�;���g���a]1�(�O�k��^�[ۑ��;�<���F�s�1^B��=�XdlI`�L���̉�����y�!�TK�ޘ�Od
���#��vy���9c��`k�v��GxB#�s[K�h�����ak=٩$�ũI�[���jx5�]��$-������р�#[�G6Ï��}�-�\r�%�bwZ/��=f@����?�;=�
ԙ����z�箺�o|����~��*��z��Σ{ҡI�h%;4�G�}0���~:M�g��%  �}��·n��F ь"��+������sڴi��,��epi��q �?�я��2�,�j}뭷�\~��PX�In��-���%�o�����s�L/:\���'�~��?���s?��f"-��}$����$�Pe��H3jV��n���ټʅ���#�=`%A۠kCX|��m[�|����ǡ�����ߧ=�� �&j��0��/]R\�g���зm��+��������s��x�v���	��/¥��k����.��:�c�n's˴�	��$�֟�����/6|W����Z��e�]��s���T��9�6q���%�ǣ��~�G FK�ː����‑9����ޑ���܀�_
���{�ӦR�$�B�O����+V�XQ@�b���'?��/~�A����9�<#��-���Kj�-��sb 8�VV�C	=H"ft�i'��ɼ�t$�==]�����{�Ԥ5�<ƁE�O�q�xJב�����?��C=8�әH&�s�v.a�m��^ǲTXp�D�dlkk�/�+�8WY�h���M��=���A�4L�rF��vt���W��� &{'rY�Պ,��dɒ_��צʵ21�w�DP��C��+_������ԁ.�pG���C=n�G�T��\,04,�w��]�,�}IK#J�bǃx.?�[4B��V`  ��}�srޝ����H�,5�� ���L	��n�i��wgG�ЖB��O�n�����Bg�ܒ7��\�pSRD+R�K�-�<�=��Zv.���ٓ��c��/��"շ�6QWST�7%��"g[e�8<s��t�AtqcNe9����ui�h�h�w�yG�=�,�������� C����zq.���>��p�B؂���-9����C.�����K�aշi]�&��K�����v��(M�/��ĳ&��+��j4�!xOFg����L��+�ܤ�n�V��f/��I%	˒e]�3������2���.������������s�~��>�Dv��倭�8p�%	D�Uܠ��<�P��r4�?��j��y��f�ԩ��M�@�02>�O{�b�F+�*��g?{�ǒ�!mж�+/��>��
�\�,K�[�n��|�q�G�ڶi�Z�ʇ��\m*Te*��U��3�---O=�df��|w�j�9s&e �
�׶�	 +��0a¢ŋ^y��_O9�tWgEUV���K���%?��Oc��7��)�������m�o������l޹z�qӟ���P֕QX��<Qԡq���Wd��[K�c3���}o޼y����G�M`����ɨ��8,���R
p'f^:��u�m��3�.`OD��H>���W&��d�K�����]+�Z��?�o��F���
KLU�Nd�����o��ϋW�ip!8+���@O�F�%� �C�c�X/ȝ(Y�nek>pE0m��o~�o���l�����H�͘�E����"�2k�ض�1	2m�3Z�$b���������<�@*�s�␔��'N��5C�[q`�(�E��@3ӧOg�^�Q3���,����?��b�6��Ŕ^^"�V3�=�E6�W��A�ab�+�\*�QjgQ��K7	x�倯��������1���ҰE�;��_@�G�������9!��.����@u�D,���`��|�#,ͤl�����"� >��,�}7�K���t}]�J^|�ŰS�L�0�s\Η�X�j�	0KΒ��[���(%`q	A}\bF�i.�䊛�|'�������k��ʞq�XH?�w<��8���W4��7����� ]]=p��X"4��=�s����Y�
^|�ʕ`X�)�G�BR*i@�AN*�9����mڼl!յ}�t�SX��s��0A��Ċ���!hXz�v��R�lq���(�5�2W����v��g?�Y�A���dr
n�����oC��E�(1>�3^.��rq=�Ð���?��K/�w�WA���ill���?L3J�+�V�.�?
++������ X X����C!��1����mȍu�v.�}�a�hx���o�F�ōSb<A��{�����?���I������뮻vꩧ��v5�Д1>��n���1���#��MMM� ��#��� kQH4����d���{�w䊜�U֘���ۯ��h�ѣGG6�ͧ�N5[jlX`*���9��Ce"�`B�$ �e��88��6d�N[�4�l�jH�2�犯j�_h5ux��tӓ�P�ysVC��\/ݶUm�VlM��i?�/��0�&M��ٝ�q�M�&S�L:�n���zu�	O;�40�)�'n[��/�Z����?���-m8b����z�gʰ�m�LdÀ�c��#X��{ErɈ�"<[	�`���d�O-{�҄���?�x���˨����Ϩ�э�h���:�����	���Y��ߙ��nL��R���D�ۃLЦ��s�7�����oQ[ݶ����>3�P����4�)O��2��7�/Z�B���_���[�6�}�gB���WQ2�M�	u�?�<�_(i�*��o�e�YA=zd9��c�O�>�I	�/p��~��_QgI
)��0`���B�0&4�Y�X�J`TԪ�e����aJl�){�3f!�-x��/�0� ��p�	7�K�o J��L��Au�6���;�<nV���<�]��q��`�A�/&�3���8�b�䟀_�����?��Z��4�#S���i��/ߖ��	��q��R��XH���@}3鼄*���S,8+{���O�6-i.�E2Ak=�SO=���.]
��t0�D�4r��m�`�������?hА�o����}�9�h��`��<�n�n�iﭩ�h���i�*m�:�'U��e�G�~C��lmR���<	%�0g���ՒiGvw���N­��
Ţk��ڝ%*���0����N��2��h��0CA,:�t���TBG��w&�7�i�&�_���>6b��I�Ǉ숂O�Hp����VŖнr���Q���b��0ӉF��n'?��\e�p;h��O~ҳ{��˘"~�^u�U ;���-�9m�:��s�Ŕ��	�}��є�,_�`��~��MŐ���l�?�[X@��c_�җ�4����n���8���ˀ��S��"���6�
�?�C�ce��|�>=�lNVy�@BW_{͚5k,���b��� J"�唗΄��\:]V]��nhh��~�	��RZc��fi�\&%�X܃*_�r�cO<�2d��ċ����O6l4�t�Ch�8��9��W��(ȂuX����&�Z�Ww�K���Vf_���.�	���P A�>
>Y�|9��(��^4p�7��b�O}�S&^��h#~�2=��@?t΄O��̟?���.�@�~��r�&Cv\1D��o���� yK�~ec��0|?��~A"I���&*Oh0���&	Q2�����B�@�/�ˠI�t�m�F�|�gpJY{'�!�=��ٳj�����an)k��s3���`Lqg�
+rR��t�����캡����իW�g@���,
bb>`�/��}�]Gu��{�ۦ�V+ɒ�U�d�]�l��ml�1�0�'	�$BB!!$T��P�)�-�WY`[��]Z������7���w_���yz�޹3gN�Ι3g>��3�8��+!�?{�����aiYH^�Z��D/�h�_��"-�����!��?�=�(��#2q%�����Es��z{w�a��؆���Q��d�p5�W��N��m�pa����ޞ>�~��}Ϟ�}�k���f��J,��v����@U���o��)��_e:��=��,Y�H�Xd�ʕ �K�.�T�?�J9�qܦk���뮻�7@!��w�V�޾>=���\b�Y{\��-pY�B�� ���4�s�� I�z�`볎?�:p� ~�ήQ�޹��X�м��i0��>���}x�܉�6y��ns6�(���}�K_z�ǯ���IsgΚ5�!�ȱ�߿�	4A��@t��?)9T�WCUc���!�[}�ѷ��-�mM��F恠e�ڋ/�c��"$��;�����2�B~�w�]u�Uo|��N�jO�vvMA�*x/z!��R��#k��7���9�.� 4'�]�$
���_���d���*;�@封��d1S�|�;��La�ze=P��1h���tV�D�b���~���&�û�1��� � ^�7���<���ƍ�px���UNl�=����~�+�#�����܆������ϟ�!w�\���k��|�͘.4S�9�mS!��ѹ��I3�B��b�P/�g΂;:o�\|�%fF:��}����A�F�.W���QOoh5g�,n��lm��(��<~�S����.��SO=N]G\xx	n�G�N�{��L�:�n�#�ꃱ?��s,X��,�K��0ѷ�r�Bjd��F%���ikt��>|?�����>t{ܸq��5V���3����I���xb��v���z�03g���|��h<�Q����2�.jux�=�`��ٳ1�$>7 J�Yh�g�y��ԝЧ�K?�k�	\1����+a��Z�X=�<�Hr
�"ylS��F�oS���>�&���kע�/�d1>��:! �m��v�]w1\��!2T<:�nꙧ�!�_r4 �M�hժU����G@����9��-f��7!�'L���������o��]t�U�����٢�}���Ý��c�?u���eֈ�vyN%: ���8묳�Ƙ2*1���$%�I�&a8�� �b6������	�vA�c6�Y{�1�ŋ�o�ޅ�0ӘX�� 8)cd�ڬ��:9"ΐJ A�,fN#T�M]��n�0�	�~8������h��ā'-Z�QH1%�i�
	�U{�B���)�X�$�Q�,`BB�BH��Y\���_y����R|�+��1�ӧOg��CC��!M�n���*�%��@����kkk�f�� ��m�~A4���BS�I.t�Ƥ�Tu|��ֺ��/��SN9E��f���At��I&gŋQ�W`��	�}��'�ۉO��=p<�[~�aXU6[��ձ����ng�.�{��x`���}��c��X�>�2.w󃓠�M�K,X��1�Y��{jRT,�-��j*�g�bx3F{��?���uG� ��\��-Iw�5� )�t,�����F�� 3j��D�&>q2�� ���`		E��C����W���'b�1&i���po��A�SN>ɞ��Zh�[�l��]; ��N���޸h��4�L�9�ZN�4s�ܮ��mL��h+����sOgOz��Wذ	n��5����z�ih��cOn]��ĳaD��Qw��㢠9��m����cO�~��M^ZѾ}{�����|��{G�������3Ϝ�6����I��v%-�g_;L�&3�b):�o~�7�tD���`"`������*CP�Hf�6�Kr4�� �x�i�A�2;ߓ��Vɫ��I����%!�K�Ѐ��0< [PRx;F�CZ��	ҍa9�cF��~1~�.ڄ�����A�0�$�:K�\�]����Ɵ��"C��z�%�$|]4�a�@:7�R� ��<���$����=|TH�J��2&*9��"+�F|��� )0�R*,�+[�ly��잢��\��X��8�4���b��6�,Q�O8a���9ɣ�>��z���.��bt����� F`���Q}���/���ij��ݿ8������0�bl�QC�0�x���n�.���0�s��gq!��I`�ԯ�K*H�3�+r���(�x���ɓᎢe7��.��;w���	PɋdF�qؓ���$_�F���&G'���˰�^In��t��Txr�ĉ 5: #^�S�ܹ�W�%��d��@;��{/%��!��MX���{��W_%���IC2��'��P!P3�o�� .K�,} �x�U�g2k��A��%�%��-s�u�� w�C���[@�8�>R{D�
n#�.��r��w�=w�0$��9t�CC.}y)F��@��|]}�/v���8V���(gwάY#�E�wO.�}烈�ׅ`*��m8�����������fN�l�����?I��Y �`�S⸂}��y��w�� P@����1�v֘hn*��^~��2�px� L��O�J�H`D�aJk���c4B�� �� V`H�1��1��FCV[A��@��	a� J`��;������a3W��L��9�<~��߿������3x5X=��ë�'
��xW*��
<R�;(p�v´��tq���=���4��/�IM��Ν�U	a�r��{�h��]6���Ϡ��ׅ �A�F�b������o0X}�!У��=�3f�'�'�J�e  �v<u��)��FUc խ�?��Ap�ԩS	]��2�9� ��P�G�h�4dz����۔Zlg�,�[�R�a���m福H�9���mF�u���=��r9e����.���^�V͸ñ����HjD5�Ȓ����3��.؃��GI�+�^�/�3MD�ڳ{��-�oр��g��+��Σ��c�u�J`s��Ol�:�*�$����F��W]1Ǩ�l�?�}�;6o:<�b�a�+}��q�l)���s,��D�ݝ���g���|�c�IޞP������+5]HL`@pXz�ΰ15���$&�Q~�D�MU*���QJ�3 �
]|	]����=W�5���ry�p����m۠� p	}d�BU��<�]p��I ����	}L�H��a=^����z�?s����Lkg�ڡ�#��u tH|V�H噾�-۔���߯�ܶ^t���@2=^� KO�$l6�{$f�_�_�z������)6�gW�����i����U����;��>~���646��P\��'-��� ���X�' w�֭Е0��uּa�ߜ�(���Ѣ��3��\SƗh
��O]fK��e�mΟG^:k�G�(n�����)�F|,R��F�T�D��� ��o4��n��s���ke^���E��w��>��J��8�@z��N��e�� �cjK�43��H��8Hn��;�$W!�d�������w������I�p��H|桘a���R�=�ԕ�#m<�5��NF%���u�ƌ�w�$>r�0� t;9<�	<��u����#��gXʂ%u�O]��1�ك�[ZZ��1}� �&͘�E<бׂ��;\�0c](���]�8�CcR�Iɜ5Y�J})!��M�-򽸵��J[V����l�|h<rM�vy��E��'5�<��}��Q��D�zQ~y3Fg��5�z.~%��_�@�V��8�LX�{��/k��Vz#��z;���>ģ��IU
�X�x@ϟ���L$n1b� �[��h��wI�����˟\�.&���$�^G������Oѣ��gw�)�SB#����/k�@��O���5YE�MZZ� s!S��K$﫯��}��pBC}3����xذ�2����fD�$_缐�bO��;.����b-9�M��M��-��L�_|#ň ��oh����u�咦|So�7��9���N������`BfQ>H֞Ii���
�_j, �&�H�R|(!��Lꊟ�xE�j�Q����b���Az����f�C�
�S<��UW�+���v�|��8jʔg�]�:zf~��4��(m�=���=�%.t�}̢��f�.Ľ<���;�2�w׮��\p⚚m�1�\��zL�sE�|.��Ҡ��p��o�����:r����*T�(jOa)-��hHѢ�HK���W��5���$��S�qI�q�� n�qB��4�\�K�P���1hJo�ԼQ��j�tUF���d-�LyW���♡�QY�� ��1f�PC�_�[�-���vK�H����[~qt�&JP�qKߌ���Wc�j) Q��dEk�fΜ�����2���}ݺ�� �KȅÛ[��N]��Ά��v47�Ӳb��;w����������]�.���V��b�W�wLU����\�Н�؁�=R%��otPk@!r��{N�g:xR�Ir:˕X�=�����}i�'e�N�̾)�j��(�СJ	|J�Q"o|�cfo'jQ�}R_�W�,J�k2T���n3�q��I����f$q�/�\�>RZwÔ.��EQ^���O�h�/[�䥦��#?�w�����Ls�	n�qY�=}�����@
۪�-���a1�<y��ɓa�7o޼qӦÇ���`�h��X���|����������(ɺ��|j���(_W,��NڈR�,<iW�N()��2�c(��4#��	�i�<�T�>}�����oL«���D���b����! rpk�,P�MFTpgiӀJ}�틺�h�\k�X�$�;zOS��R~%~1JB6F�6�^�3m8Y}���:y]���3� 6H�ɛ�JfƯXJl���4R��gn�8�gjċ�Z���o��:3�QQv9f4���AaA,J��^=S\^cUA�HeϤ�Y
�����a�S9%������! w�V�t�Rҝ��H�n �Pk�������B|(_�z��sa.N
�婣��ZH0���$$,���@A��2q͜*���F��ŷ/r5F�a��������O_x��'�p��1-xK}�؏�+��Z��{���̙�Ѝ/�О�x�0�lGώ}��X�ڮ͛[�1C
�q�W7i�e�4ܷv��W�o�i��ΕjC F�e���M��q��O��J?4-��I�/F�����2G��t@Z����$�/1?BְC�xݬVIl���1�5e8�u$4t3^x�'	�}S��?��ġ��L
��QV��D�x�-�z��'N4&�[2��l�V���;E��e��%Y��ql���&�x���#�o�W;�z��a��#GΚ5��rcǎ=���W^ٶm[�r�џ�-v_)��n�ͅp��u[r4��x�۪X���=Inڸ������uژ"�M�	�8���)	oD����|�	�e︈C���{B�h�?�|P	�e�u��O7׮�@�������gDR���2�/�L�3����~.�\�6�K}N�4(��xA3ʟ�����^Ο���9�p��R�Wľ�Y��&���j�έ�s!����;����iՠ����#�[G_��G'v�n��X�N��"����9��cƌ=�S&Mj��)�.\8��eٲe��:�+�
�˞6��.�o^��nޭ�ٺ���L���6�M�f͚�;��ڵ���[�DGst��"�|-΂/<�.��*Z��q��Zd��/ĥ~�u���3*6�4Gp���?WZ�ɰ\���#���b#��FQ׵-����_����*�IPT5 )��Xj���-E_�S�,��(���/�H�L@��[1@ƟW�y���rwH%���k%/&[�r�?5��{����H���_�*������ԘJ��)��Bݦ7�\�'B3�܅�iy����{�#�QcK��F�B'9#�I�#@�DJ�qvؿ`*��e[��?�~�`"���
4(-]�K>��A�Ѻ�\�Ԃz��Mi1JiM�N������bZ&M�r������G�����7���}�a�vv?��i;�y'��S=u�����a��/��qX7m��%�ׅvgLG�<;�HOc1���k��ý�q}�n�j��S�ð��a�m������N1N�&;-z�%z�Ð�{F�$� L}%��F�)�_�b:�����gAA�w���ک�W�K#�E���҇�i���t#Ci_\�LE�3t��:13�(��X�o9檅�2��IYڥֶ�Z��M�1s�v�}P���q���̝�E��0�Æ?���n��V�(�@$��a��7n۶�4@?n>e�IpW��'���`A��)�A�&���42��1B:fJ�&��efJfP��d*�8�@�]_iS��+ʦ�J��Q�k��)��1��u9	b�1�� :�����d��/���/m/2W�C�&L�Dh�+gH3��Y�8jS�Z2���L��2��<%����m���*u���y��L�5��̓�1���;�Eu�]0�4iJWW���������sv��^��r��;�ؿ���>4��g.���su?�pw�� Đc{x������H��Bf8Z�D��>�D�,̓��;���c�[� p�I:�҇c*I�~3�-�4����d	^J��v����n�K����:�n�N�7�:�F�V�I�HX._/Z-��L��M=�Z"��4�6J�f��e
}�7+'x������yP�v�X>���p�V\�P� x����2�&rPZ�!M��5k��7��m�_�\ll#9YQ�|��رܐs��0���������ǀ�z��J%�%rk�J�K�>�4�{t�f��C����}��a]���Ӧ�9�đ#Gnض�9$k׮�[��7\�7n��d[,���oY`+��>�֫q'D�X��D�Q�����&��9tн��)� eD��{� 4z
P�v>��u�ԭ�:O*Â� ����������� ?�>;|�Rn��x	���z���%� -��ys�ܳ��7*���n��y�����L��l^�%C� �F;����#,X0u�`z���f?p� �e�d$���޽�~	�@о�vk��}Q.�P_����<xp׮]uup�A�Pl%���+��4��<�Q��2X��H¨d�!s���g�ֆܲ�̦#d�4����՗2�����H��F!O阙�!ȩ�X=�l�hC�S��|w���S�Ν;y��}���6�Fv��yi5ƭ��ϟ?��mذa��ɍ�����_^�}�v@�{�Eߜ9sƏo�v�]gAȍ�G����eR�>2^�&{��{��S��ϯH�ҕz� c�dt�20���J����8�KRg�/������.�L�P �؃]E7e�N�+�Y��+0_�҈TX����/�-�4X%`��k�T����7��@���)墠$�^�u�N�zi��4�#�ę��;!<h۲ǂ���۴~�o�pZr�I�����M 2��������|;�Ea͎:�4*�~QO�C�捷�l��-󭛤�/]��4,@��3_n�q�F�vuuM�:�d�3��z2iS��zxjCo��>k�/m(n\��-Z�kT��. ޱ~���8�79��4t8ҹc��m��[�lٿ{���69�T�8�\x�HS`�?��ָ"7&V��M��I��2��EYr���"��E��_"Bi�XÍ>f�b�E�����v|���X��U��N����2��،�4&׏���|�ՠש ����L�eJӨx�F���[T�������}`���~��ʪ�L�={6~�1c�ƍ�}}�^{��.����j=���ݝ�F�`x���ݷ���C����
�^PW�P#�u�{.�Q�q���)�^`:�N�凡Asm	���4�xLHT�'�+ʻ��0�\�,e�e�Fs,������GD��Xp˝�9V���A��������h]4�!x���N��DFs�G�8�q������X�Z�n��W��QǍ?묳�u9��	sg۴�΃;�o�:mVsӰ�N>uҔi��mi�Q���i�B[y��������c�mA���ħ�4�x#��)��
��*_p�%Z]�|�o)���k�q�~���o:L��T ��mP�ziTR��[2��_��3\-��[��~Eo�W&,h�g4bܨ�%VU���s*a<�`Bi��l��*s_�h�	�;:���%6�o�o��t.����O
7����xkZ��c��>��R��3Yt>��ID�7ր,��/Y��X�x�`��;�`�ԩ���ڴfh�a딍5lԨQx�ܹs_~i+T�+��2cƌIc[[���N�s��}޸qcgg�����߼�t�Y����*u�Ses�{���y[��bz�}
"GU�5<f�xE�v����/3��|�CԶ~#�0>�n!���x��G��p��B.�� ���mf�?�>�v�3q���~��	|��W���ʩ\���8z��.v�D{b1$��m� {��͒{�e˖Y�f��a�&N��~�ܹi�&��X`��LY�*d�_�b���q�z���ZE萁���VUFK��u
�P8q��2�'fHQa2��d]�|z��{��S��ҝy�)�n�^�Y�5�K�>	n�"�����̱�z��#*���?�4#ݔ�9r�i���&�lվ�.^��]������I�&AL ,K�.>bo8ϐ��S�#�[�z���&wŶ�D��>�0��8b�~����2�)��5��T�t�P�H(l�����:���f">��R�B����5iR�'ܒ��<��z�w�ƌ��� ��/G:���=9�X�s�+���FE�̟��m*������C�lA�n7�bN3g�Z�I砪���(Y����S���X_�����[�M��Gw�������g�*�w�h��j�o���>�/�J��QN�������8M�2h��]ҁD�Ɨ�5"�����R7��+��̰�V�4n�vE������۶o.)vwF�-i���V��Ҳnoׂ����F���3vN۪5��-+��i����?�wڴq&������lڴg���G��A.f��iOo>4Iz���
4���u��Hc�oɘ��p}�����+�X�@�@�O麁tkT��lUg��V١۳H���2���Xz�8b�C�鐢,�/��5�����zyF�K�2�|�%�h�c�~�veb���[Ї����/в����I��Q�6m�<m�T�,�b�W�4��۱�����g�nL�+����yh���ht!�u�{:ѱ5��ݺukב#9W�8����W��/��	Fe������y������.�c�L:����������`�˷2G�p:و��C�����|tiiT�ɍ�	3��Mڿ��T�"IEҵǥq�J��%��8;B�(��W�:���ճ{��0B.2��e���X�r���N��S�Nܼ~C|��O<qꌹ�;�����#� G{vo_�a��z��]8s�����5O�~
ˉCH�I���;h>�*B^S)��O�uL�p�Lw⳱k��:����g���-u�Pf�=�P૥�����Y63@��b�
Lm�U��x˦TBeCՉ�J�MF����%�.P���S��^���3�Ӫ���*��`��
�����i`r---p�[x��؍��y7��h7_p�m��B�$������*�PS�}I���@�L�G�a'�z���3*�{LQ4����3uZ�\BO�Bp�w��n͚5���cƌ�2a�{4�;d�gT��ݻ��w/T�4�X�֭+�]�.>҇o�5+<�\l�{L]d���v��,=�����=�;��
���j1��hh�g�Ko0�#Bm9%R'c�iHi�F��w_�8F��3a��WP)% Gϰt�vD�"�Vd�U�)�R8�*��J��Վ�����X�̩.��[dX���(�6��R1�[7o޶m�ȸ�f?�u���+W�S�r�������ڵ�7.�[�nw�[���r���ޞ���i�Q�*���s�ꚩ��CDF��4�B�Tm�T����"����[�L�.ʬȑ��C�S����CjcLFZ���&�#z�:l��3�K�{*UJ��˕�V���V�?aWW�2j_�[R�4�/_>i���h�ر;ڭ݁�/�� ��SNٴn}1Nr���G��X!=���n���߸:2�I���[r��`]����]�Y�g�O�1���&_'�?��紲x�� �O:#�;f��
Khg@pQ�O���0��e�����)!y�B!��?��Q��BiI���h:�8#	���Y �h�!$�������/4�	���CGXLY.t�)��%l�~���8�q�ܒMSF����us�X�G����V�����U�:��n�&�$N+�+d�E��?���H ��F����pH��FqĴ`�PsÆc���3q��H�'��c���*;��B>565^��V�책S[n�/��-���Ў���y�vnٜ6vm��Z��v��?{ܴ�c&�ڻۦN^�esC!N^xm´i�uuH�E]��uL˘Ȟ��Ӕ3�q�'�z�	l�δ;�[�s���C��������9w�B�=����� Y0}dAQ:�I��zS_I��	�j K.���4F�R�����-�������?�m�.�~�]V�⠴�`/��Il����3XO3-�o=��Ũ�-�݅W9r�:����Qh夨��Acˬ���<4�;ڍ9�a� ipW�
"���b �=g�bŊQ�F߃n������)S� cΙ=s����˂�<|��{Y�}��������mz�
.Hi$-�*�K�5�� �#�6� K8��z�bfļջ=��'R	W�� ���e(.�ʡ�f'CZ��1<Y:Ckv��tyN�>�gP�~��s�`D���싲K���_��D2�'p���!�����S,J�m�Y��#��}�����4�� r��;�B�3z7;w�3fLS�k�I+֮��^��г6,X��c�:u��o��Y�P?���w�mQ��iW�[���@������@�VP���S�ZZZ���s3cWm]t�FX#=zt�+S��`H{�2c��,��sQ0�Н
�#Qp�#�����&��NQ�H������i�\Z=�$=vj�6��>�]r&�k����Ɓ_��E6<��d��u���]�:zh���Y!���:3(��.Bv|I7f����0���-����s-j/2�'x�	K4�h?uu�V�Yl`Țw��ǎ������.\h	w$>x�`�����u�s�L}X�E>E��tK�kD���	&�z�g�y�����I��={����O?��ڵk�C�Azo�OD�;w�g�u��ֆقS�Ɵ���K�n۶M���t=��J���~����ds������W�~��_x��$��Q�M� 5��6�m����={��ƍ�d[M��"oܵ����g��=;w�#��Ɏmj�袋N<� �Im1y�;v�^���?,���/.��?��U�	cs�8o�n�0�������SN9����P�nܸ��_\�lh�9Hr �l�Bk ���;o�<�3��M�6-s�;�1l���fkk+���Ϟ6m��b6W�Z��sϭ\iIL��?�q�ԩS�8f�C`�k���c*�m4^�?>�_�!Pa|kҤI^��(��<�����C�C��D>c����O>���yV�-[0�/���dT�"��$L�����8��;� ��a6~���PeH�`f-Zt�9�86���-��g����`UR�۷����O8䲈,W� �������~&X��b�S�6}��%KN:�����#�����?�m�v;��2g���ډ�R�v�i�	� �M����d���
}�k|�H!J 4h���m�?h� ���Q�_098Z��K��ل*Ї���109��w�!�;�8L��^�d�[�jm�`.�{p�[f͚Q�Xm�n�ڴ	�HU�9�q ��.|-4�ơ��Th�_�f�*}��ݩ?��Y��O<�ĳ�:kΜ9���"Bf��g��+���h,Zt�-���1]��t��)�b���˹���X^�5 � ����볦����<pš.w�Q��rʩ����1��9�ܾw/��C�=�W�l�_ԜRb�
a%�7���ŋ'N��^�&����zj���O�<L;�v�<I�`�
F����L~��0
�ܺu+���~xǎP��ʽ��dv+FQ����.�q�T^1(9��J�����AWa�@y4n5�с��2��CI��aX!D�c��p���E�ɠq�NM�����*g.�w<
 �BJ�QB�hJr׮]�JU��\P/h�>e�,�"c6�x�	���^�P��;a�����$�/� ����ի׺;U����Ң=g����[����'�Ҿ��muI�\؋o:��F��vv
����[��$�gF>|�PC�)�(əB�xtw:���I�6�w�t��r�W����!`8�w�0�HX�������z+�D�S�Bu�LX�Ͼ�d!|?{������hS���|,*�����������Ye}�!O0�5�\��w��Ε$��'��<�����w_z���}�w�C��&N۽�^F�jM�	w7Duc&�5�7��?:l:���E��������L�􎌷��<���7�����5�A���D����4,�Æ�Imm�]vه?�a����-װr��~��_��נ��Y��V}��ދ{���]�B����Zv	��r�-�>�(fVN��y̩�z�B[����-oy�;�	�Z�8��6��#�<���bIp#�7z�zA�+x��xz~�y�q�Bp�q�_��_�L(Ү�(^R�(�٫�?���E�vf ;�J���\���/��N�=Qza:-MK͌��h<	���D�+��� �����;���{��P6���S�����=W_}5�O�3��>Z�*������~/Z�Ҵdf��j+0�W\�$X1��4G�����瞛n�	o��ؾu��	x׽>�3���C��i�5k䬽7��~p��>rT����������V�m�������O�����7����"��6�x�����X~�C�������z�b�����3�@����ψ^������.\_|��^K�3�I�͛7�{��6T��?�ý%Ǯ	�C�W��P��r%as�&���OqJt�.����t	���Z������\#�������'?�	4ú�j, �P���. ���o��B�qK�(Xh��v؎�{�JrZF��s�8:N� {�| �!�J����|���6O=�o�i?�!*�R:z���~7�>&�+l�a�����W��̿ƅ�-�:�M!d�mo{h=���8|� �o���={�����{����0Ḱ�^1~h�qO/�e���&@V��*����2�5��c�D	^̙�;V�>0(���dp�]�h��/�������@�s�͵k�b6�����u��6�|��r��ozӛ�� �,��Jt�	4 ��	��3�H�:Q8s����ѣG���g�����Vv7@�0���v��ի%*Z�q�RR�i~�p�}�\̔lG!�@��BA�C!@�03J�>�p|�� [��M�Op�0�0�@�<�Z��5��N/��W�,�h�=���"���0 �#�)�������B�,�c+��/: :��w�YiS�B��z����P/�6����m���ɀg�dx0��X"&�j�������_=�"��8�EV���w�u�N�t�b�!�y�Z�����P�|�� �&	�i�&R��VH�v֦L<��4�\AH�ECd��5���#�����r�ǾI���_����s��v3 �w¼��ͧ�����xݕ<h7fuɒ%���7�w�*�����k̿$������=�������� ξ�KN=��0��_������%�+r��>�я��_��	'����F��Z �m��7���,S�N}��?�bjK�\s���K�W�l��\__c��O��u�]7n�(S�8X?�5�����68����x�b�"3�S`����=f��ݴ]_��ñA(0���4�o��opʹ#��N/��`CT`恇�>�!�r��,L)L2����E�˹�������ã�IfZ����o�����D2,����&xʲn>�I���}m܊�l�D��@������`��ʫ���&YĬ��?�P(F�e��E*q��s饗~��_%��ebS�ʠ�?���8��΋�pr\���5�5�f��(�)�C�Os�>x�aZ���0eFEԈ�'O�ҁ�7�pÏ~�#����1��7��,�4�0�5���B3|�S�� � )BN�ϟ�Lx8PgL$õf���}��ouf͚��/~��B6{"�z�q�����+���ùЇ"g4�to�U���>�Wp*�ä�ŗ���s�������������t��҃{�7�!�7�p,�եaL��'?	�C�N@�Oq%$>����~��o~󛡣(k�������K������o�D��r�*^�~�cځmL��`l" g��!�eg���*���p�E�+�,�2o�c�F�j� �A�B��+p�k��@��+l0��>�3�����0�5b ����̂�:h��'N��kͷ��e� ����/��r�-|�	eN��8@ѡ��C=$�V�Џ20 �n3d�������.�}�7Ϯ�~�K���iӦ	mc1jt}�p� M>���x/������2�A�8� ��Ip<Nf�aO	醹^\hx�\�Ԩ��3g�;��?���7�hJ�ä��Q���@������?3dR���n�t�@�������NN9�y)�l���!�i�Bf?���C�R�b!!!nJ���ۿ�[�0h$��P�[�}�x��?��?C�`	��#F���6�7o��.�iV�F�&�S��I�%����d������g2��ų����;mmm�g��e���)t;�V�q8�쳿��oP��ǪĐ�m���$`.�Cc�1E� h�{�Ǿ����j�	f�_�Ҿ�{����4�Nx3�M�1�������c_,�"�u��?HJFm���G>���7�"u��`�A�������5����x�������wɈF"+�u��>y��'���e�յҗk�K�SLM�q��;
rŴ��ސ�t)*��
�}Q���L.�ˊ�o%1���\�|}]�����������uz�hLQ	A����U����j'�0�|�G��A��S�5��><�|�G�>Z��W�T_����Շ���㌕F��i���|���n�	]6��/~�Gzwu�|�ىsf<��sf�~��06Ÿ/
�/��?A�s����%qT\����\�s�X�f��|">|xP��o���3�Փ8
()X � ."���|�щ��@B�6�Z�����5���`}�����ﰚ�6�y�/	�� :P"�Yv�n������@�,�=eT1-<�E��!/ݎՎU��8��tH����F�L�Qٱ?HN����/�����o�3�iE`�X*(;
4�{7�낞`����K/�3�{��<�e�x{z��K�n�P���}������x}T<�EO0�qi-a-7)�41�/~����J ���N G���Ç��C�������sK�Z��6���҄(��^~��!�,
�,�j�݅�À���-#cۡ�bH���4��p���%5Yx?`�7�������':<)�C3&`/����ÖӸ%��/��o@�T��X�ti���՜^^���F�7N��Au#d�����k�H���y#u�ФJ���k`E�^����n'd�����p��s<K�&e|D�;&�=�7j�SvO��`v�'K �|��/T��k`��=��O�ӫ0�`S:up�� ��ғK47��$(8|x��y�V��O:$�?�g��4ܻw/A-��?0:��h2^�Q�����=�\�ڈ~B�����0)x�̣��> ����C�W˃����7�pƛy��6hp������c�o8��j|��Q�\̗Hh�� �?�ǃ����}��&1�<��a��p�B�������&4tH�k�����W�ZE馞1
��~-��<�>8}��#M����ău�U�7��y��_��n�#0ܒ.=��?���ŋa��뭷��%�bi��b� � ��
�Dͩ"����ꫯچF]�b�A�w��>tp)dP��ǡ�\��u�]�a~��g�A ���$�F��S�HP���M��Lh=_�`���i��U��G�,x�p>)DriG��6�n|��3q�~ߴi�%n��ס�Bo�~n�e��$��j�)UUf�~�n�� 2>�#A�����0����`�׿�uh۵k׆���^]��b��3g~�K_�={6=T	k�3^���o߾��3U.��7�'Л��b6�*`�͕!ï��y�5��˗/ǃ���(�����3
�Q�{뢺O�3�x�;
1�{��&��Kh�\��`�_���8��P{��A2.J������m��W�Bfv����/|Ar�5
)��4
�����Nn}
8#�4P�����#�"l|�\�q�ˤ���	�d&?��,���=>�f�i�Ԋ�ʰ�$0�'�� (	�,0��Wc�P�ݝ;w���r	� ���E�v�,��|&X��1�B�� �p�2.��S�.X���SOM|�&m[�+�D�~���$�կ~f^L�Qi��F?��мd���\�q��{	�(����Dg�^��ys�*�h"@���2g�����ɶm��������d!n��9�]ĸ`� w\!�SUx'�-�P]z�`h|��Ie�ȥ�e�8p��idf��{���z����Æ0��	uN��[�K����M�b�|DcL��Z�+�l>��3�_|��2�=��0@�~�2�*fSp��&D��v9�%�j-��. ^v�%~�,�|���ǰ�4H�YN����g�A��p�|�N�H�����rFc_B[�1����{ ��� F���Ǎ�n˖-7�x�@M��q]V�SM�W�U�+���h+�<h��K/�I
�Y�?!���g.���ծ�6M7�~֢�!��#j��~�s{;�.[�~,s�W_�������,�&q�v���M��M�����%��'�$�v�v��%,����?g̘E�لGĩ7^k�����{/��2H4�Zu�N�^B��z4�����4���'�
��}�`ڒb����E ��.�������Y�~Г�$i�Z?p�.��r���R�
���f���dq���"Z�/r2.>@�_��W�ϵUϵbt���>�nZŨ�C2�4a�$t�ƍ�DVZÈ���Y����O�	J}�x&�I�}�O�	M��&'ՙ� �����aLEHId���2��D
Q�^���D�����..T�hJ�M�>�q$���/�[���G�a��I�R�r`�
fh--��R�a�O�1�;ゲ����\��OsiW�=嫯�fD�n��q��B�h����/6�0J�|c$ih�g$�;��֟�Ľ�7]r����J䷫3",�p��I'�'=6���"�f���s�9'p+ș�TQ%�'Y����w���?_���ہ��c���"�]�L!8��?�����=[6�ݽ o�Uhln��>b+2��M�>���~�𖮞�Ɔ��z��Ή��lJ]��#�t�����lq��+�`��G�K��-�T4�Ԇ(���?u����\�S�J㝊�'�~�5�;����^�:*M`��R0v�4N$�UB�[�S<h��)�17Q�[Ȓ����w��~3���5�~�X-�����p�����+��'<.���HB
Y��(�*`+`1�#��3�2�o�op]`�R_1�������.����=���?�ꊂ�R��gAv�	�,���5�2⌳{ �pr�z�)�r��C��.\x��ң��/�t��<	��9|��O���}���_ܱcGGGG�����E3, )�%���ӹj	}衇n���B�����V���&�����O�?�V=���Y�@g���W/]�@3F��4�ȥ<���ϟ�OeRu���Dz��h�OH(��x��F�E
�N��h�3U.n��B�,Kⳡd ���K�>	,(sg�
��	����wA�8L�`�OA6^󰇐����'��뮻$I:R��E_���(�C	9_�C�� KLM)��s���)
�^I1EkP�%Q���'OχZN�� ˃" Fyt� ]���H˦ߝ.�Z�h ��[@��{��ٹs'  �g��K���ژjQ2*��g���s�=W��B� n����æ��HDO�{�LW��'3��]�B¦��>.:`�|�O>���_}�U�aˣ��͉d��o�G��qU0�H��BI�'��(?ű_u�U��63[�Ԃ�E�qmrt��w?���9���&a�`���qI���MSƎXn߰a��w�\
d	+ ���PF-�K�e�fΜ9@2�������2�@2L#��H�Q��3�_q?��O�����˹z8�	��T��k����+Qݩ��A��E�pC��L��[����Ap�����g����p����G�[�o�^�O���:�,p_$B����:E���7^��_��Wtk�*�Xi�7vÆ�=�Ԕ�n�w�F6���U�˸E�i!쀣~��7�:��(��-ï���������Y�"&�Ud�L��� �7�x#T��2a#.��0��ԯ�R��&��S}0�s0�r��}��U$1������{g�==:��n�0L�
d
=�淾��ΞNܚ�	��#G���`��Pj�l2t���R�$Z,��h����+��*��{!F'<!1`*8�}����ѣGC�@��<������jCَ,�ӕd�	@i,�F'����k��V�.�.0i,H|Zd��j˼�NF�q�_���3τmKTҹ��r��k"vD��n�hE�Ae�@�#��7��&��\�48�FN"C��f��dQ�q�W��	_R��*���P( �,�J�	ɢ��Di����| QV��=��kJpɒ%�m�H��k�00׎�� s�/c�!���&���R��$���7L�� ��~��ɹ馛���B=�d�X\f�a܌���%L��OơC�d<w"c�}�ԆS!!.j������c`�!#���
�^��n@"�͛���|\��[LoS6�qZ��z��`}�RFn�<���+q�E`��ܔ\�Z��{�w�]����XQ�iP~at0BP�z��<�����cn����?�!sO�RbZx�� ��zu��:r��>��AX8�<�S���W�=s���\K����F����͚5�Mozۉ��G!/����\H�=q	���/���+�E?,_�ܨ��T-����뮻N��s�!���R�0�a������{ｷ�}��O?MC	�|J]2��x�P�-U����A�n �_p�����f� 袩��d|���$J�/<?dA���(m5R����
��G�wi�e��x}A)��w��l�pZ�!AI��K/�d�XӬH�-P�,�Z��Xx��j��-��2R�tp��9n��֬�^׉JKר��&Rԯ�.�Z���|U9}�t�����6-��G%�� >4$�����&0Fl����e���w��I���v5>�q�v�F�7ꄾ���@�T;ԥ�$п��I��~e�� ���@���@[��V�n����/Pͦe�Pq9���O$�%s�ک,��DsGE��s��L�ر�CR����o��-��a�D&M�r��_�^��T���]�l���b��1�ڧ���ݎ:����8��.�tlo=��􎊊 ���Į9�(�-�e�O��h��q��Շ�zbx�9$4��uʔ)�/���R����	�chVeN���9~#���V�q���7�A�e�C�@j���2���4�=.� ����v2>آ������#�	s����_t��|��6�ئ��B~��7l��� Z�	�.�e�q��L9���*)��w��Y0+�moo�)T�3 ""i�C�����8l�����}p�Q�\ ,��."�����J\^�3lfZH���	@�h{���H����cO�G'�����0ܜ�T���E�g8�`�:~�n�jIv �	6�v���;��Z�p3� :C�&~co���K�B���h�Q����,DSЃ����W1JHE�d�G�x�y���g?��GQ+���m��.y_�$��ݸX���=l�@��q�3f�,�nx���ט����.4X:���K�M��m���u�-��7��E-}������]��$���+؋#�#��pZ0��BÙ3g���Rr� <a{�F�F���ALXD@D�T�D��O�v-�"-�k0�iܡJH��1��y뭷J�����QC���(��e����3�r�]q�g�q��?.�¨Q��2xP����ԥ��=��e��g��0#)b�c_/�&O�����h��Kk�ۄ�
��������h���j�&!�4���ru�'����3�-X0��wp��FA�`H,�ƥ��\�_Dը,GZI|��>L�4x,������;�>���4�X5?�h�8�[0
������z>�C�ɓZ	�~��A�;��sC &���>�SEG���<%�s���_��Z�=���H?���J�@��@F�n�s���x�|%���[��j��S]�{/����U"���J�>x̾�DNi�Ďh��0���믿N�G�����g�)���bV��)�2�p�qv�V`�?��������X�n��^9)"�dMl�����N:	&i�"<`�����c�R�@uJ�/��5"(��}�c�=��,��_%4N瓮W�	3��,j|� >Y�j��u�:::����N��j���ҧ���*��h��7���D���+=L ,T.w4T�Ö�����E�/4�=���l�ğv&�n�(�I�h�h�XmN'ہp$mŊ��"	0<���#0u�Cֆ��Q��>*��w����]I��z(�������p�S���O�&ďl�P0�c��_��n�O9��<P9�m��٬��|>���)2q�'��}y��g��|�Gt����ڞ�����>�Mb��_�M���˗K,a2�c�5Av�3�ם�6PT����p�ʀ
�>��v�܌s,�G�	K}�0!�y���W�@��_�*�OZ��*�*�kܬ�x�wLK�<�/#7:_��J�v\H��ڵ����� ��/��c�@ى�wɋ�`���5e)U����C��h�"X���
,.��/ER���(���!�sb��5N�Λ7O�bh�~�Z��N�?���SN/U�Se\�D�d���\H!"
[��VQ����n'������P��?"\�ȅQ��bΉ��?�x.l&jgK��7P/���b�`tIm7~f�ɇn�{n� n�2� �ϣ��s-���G�5���0�J(���>��
�'���Ȣt��0�YTeC�K�@����dfѫ:C�K$ ���X@�*��>h���p�C_�G�ϵ8aHI��^z :��^z��\�f�"0�X@Um��ҕX���g`+�!�2ř�o�|
��(��*�$U�-h43/]���`�!�yw��F8�"������ �����ũ�gX.1��C�`J5��:W��ձ��E���H�n1#�F^�$lɆ����[��w��}�٬��S�'2�@��#��� oS�{���<���\&W�0"{`�e˖I�5T���,�ʨU5�����[h<���]��'JNs҃�;ę�Y#[
"7^�����:P�\�VG� �Ϙz.�g�\��D��T��`�C���sbb8Xp,���=��ԯh�H�[ ������rēH����1X�����tX�\KnoGak[�i9rh��67&�c!]��sƆ�{l8��sX�P�	�&&)�c�#�I1�9������V2a��u����V��ʒ�&��#��xm��%T#�HG�/JV��q�Y�s�ƌ�#�b�����-�4R	ڵ�oQ��K�,r�g��v�"��͈֑�M������|����2�����ܢc��5U�O����h��+!p���&y_h2�5�G�2�	�iޤ�za��A�9�E�ѲLU��XL���h�� �1x��xH���Fa��4��hV����hb�]d��&;!k���j!�_�qe�39w����c�#Wl
�L�N���:�ZvKhR��=M}]p;h(^���WS�/pgϞ=��z1$���CQJ��r!�Gt��l˰a�\,�A^婼���,AQ�
�C�@�,&+.-�n�ߒs�4�O)�����E?K΄�sS���~֎g�i� �Cr�R���0�F�'T�0�j'"U�� �?Byq�3:�(�i	���գ�0TZ��w��U�4p�F�Ҁ�/20����)[� )�Q0Ǥ����Y~ �����X���\�G.��~I�E@(�1.���[�n�N`�PD��(�C���&��"+�|�Y	��K�X�Y3�j�����N �щ�ۤe
,s>��NS�^2D�(�
�2U��kv��)�>ϼ%T۴�|A���DA��*)�T��备25������Hdm.�/��{�W`�%�@�U���!��|턊hq��$�Ps��GQb�����ah�6ԅ,e�o1����AVCҡ@�K 3�9x-��@m�o���gs�~͖K�<Z�x������$�`� ���#���h�}BS����W�M�q=L�	������ �w�W/�����	6����<"뺦Ԅe�������{r���,���v��� ���|@�o/�&w��	���M?3I2Nb���p3��
�JUi� d�X��c��p`�9�*W�W x'��
�
�.UF��ˌ�җ�ޥ�Z��S����2�\��>��]�7�$__k[��Bšo��
���k]��޵���>�N����j�
��k���$���;�Ra(�,.�fT���O_gHWe����g�" �y|�칩ظQ�1.t���b��9U�Jߣ!�D�a���(�,�U�xy�����/���D0^����Ĭ6^���-��,y�~���8���j@I!�,���8w���l�a���־�D���dT|*T1l�[�>��j3��WǙ��B� �X&H������)���;�I�(��iG�@:�(��*rT�������;��O�Eo�(�$�H���� ���j�:���\E7����F<���	�n�)��x�b�ĩ&��語>�sÄ����-`Zi䈀j-�n�<� ���ă��,,�Ұ������N�j=�)�=����6n!���JPÈ@�M�dH誚�g��ּ:����'`ڊ�7s��m�Z�j����ql�������\�S�J%�hBU!�v�*^c��*����V*��>�����˾��*3����3�ܵT����1>��|`�I�+�h���0X5��ߊ��̱�p�h����U#5a�K�N3�����@2(e�+��הR)��Н3�����|$�/��u��5����S��l��46�
i�vX�R���ULO_o�X8:*[u����յ�	�L� {t�m��s��r�����|�����>5��\xVCͬh����r �~���y��/?t������[���إ ��z��]]�Z�Ҥ�X���Q�0�����y~�o߾�/��JU�!Zfp%����%<ue�vʊ`Ī>F�9�y��������5�g�M��ȸ�J�;�{��D�8~ŸR�UC9d�e]mC��L���P����D���_�NX�-[�HƼQ�F��bx4�J�2��:���bU�xw�O�߿��VrՏ���� �b����`�v�8
U�Y��N/��j��v��!5�sj�y�KC
��;F*�)>��C�s��5η�mv�ލ!�Ԩi�A�+F�#U� ?h7���i�iT,����1e�!�$~Q^6��ڻw�0If���hbs�P�ڗ�a����?;�ܘ��@�1Q)�������mOd���J_�NO^ψ�fx$zj&paryFM��j��~�>�}��ZT�+d��b�����S9�
:�ę��ai:�gt'�����M\�Q�^-�o܉��2�#)�5B���A�Z;ϙ;�8�a�ȑ� ������ېqGkd�Av�kܸqF��Z��Ч{|�e�~hEeɨF8:2p��L����/�� ZG?k�~�]��������7ȱ�F�ͱBx����]�3�>�@x�.PˆreZ}�H��&�g4�&8v�� �P��g�g�R[��Ѩ!�.�����ȝ.��A�ԯ��}b���%>#WZֳ�b��W��4����h�6�銎n�����c�C��9\�bFJ�׳D�K����̮]�쎄�K�3��(ֈ�G>��/_.��3*�଍�DBt$�"��+e1�͛7WT%�6�	��Ȱ�L�Ё�>wf5Fm՜�u��vf�Ν�¶��b���|uU�/ӌ�h}����y���v͚5�2��eEG_�7oܸQ쟤BS����\ n�^k�I-j�������:�h	D�2e��!s%��"۠�T��-2w���>�V��S+�ZFa�O�!W�Y����(�"֖��j������i0T�Ɋ+WlG�[�!�g��czB���A�@��,��
�nn�?_y���J�d�0��|���}Ej'�ai��y�ט��S��iC��EwA�Sʸ�"��Q�C�x���ĳƗ�6�9L\�(�n�+��"��Á��+!g�+� �D��p�nh�/�������Bmj�tؒ�:���� M���:�n$#�p�U�4�j]W΢�s���̄���}gݺu�/[#͆j��(�"_B�e�D�,�-fh��U���By����W_�3j�iA����K�4ַ{�\��"O�H2�3�����R��Һ28!(]��X]P��Vk��Ƒ�q<��I�1&�p�%��x�[�}��,�z<T��94��aޔ�jđ� 
�ʕ+k����ڵk�m%r�Y%.��FΨM���ZT@��Z�(;_1^I>�؇�������	&��Um,F
5��6�sMiѼ?���i��K#����`�q�	�|ӦM��ԧ�ӠP���WN^~A7�4I�B�n��32g�N�1C�:]���Y(��U(.�N�;ӵ�ic5�L���/iJ�B��8ivn@]1.ֻ����뱋�8��m�����Ս��BO_��L;xa��!�+l�y禶P6kP�IV���?�y��u�&�Q���=�����ʵ�j�>�y�Rb@�*ޟ�l������b��ځB��<mYAI�O̷�l޶eͺymS-〥��0	�Д̢H~��^Сw�y��閫܃�����ڸ�Z��k�"	t�0�1zN��3�|�#)�SuDP�5�7>XB%�y�c&ZI+���x�W-ZTT5��H@�o�xꩧ���Bk��/pȲd�.(��p��4D�<����t���D���0�E_�?.�"jJ�"�EĐ��-�#�9T!�¨Q��-�b��J*fAe�I�����o}+uJ���d,̥ƬI�����)>��M�M�Ɓ԰g���$>D���n�_��0��v֕�k���Tl�X�h������� g�$����4u�,��%�jtj1�		��~��G+�5uS�W0\��O0-D�ɸ	� DB�RU�R[)�2&k ���s�L��U5��������q�c]�=~�G�_���l�
�,]���n�l#�՗�x( �n}�2 C� ��_x�k�����L%'�������s��%�\�^������'�|rF���q>��@�{�G�<��:��EPes�έr�d�߉���X��rKQ��?�8π3j��Tғ����@L؎r����/�v�i�ߦ���˯���M�+���<�T��`�6�3d�+�m��gݺ{f�۬k�8��Т�����׀�-�㣏>�9��~�G����Ḯ�y
P*6fz����_|��}/w��5)��!B�F����M����A�zꩩ�a���5�_�w�qG��L�����2_�ߋ���Ҥ2$�+���,�c�`_�6�cbʄT֝�E3dtk�I�:�B���ŋ���*�F*0 �b����PA]t�$���ω?؋��F�\٩^�˅�/�nK��?�v9,X�7�R�������FW�n�΍�
�6a�����:���a��h�m?��'��9��xb6i�$N<����#%P�D���z���o����~����V=����q޼y�+N�
�,�m(�����[�*�<w�-������=8
+�-/�Ҿlٲ�{,�;��ҵ��[�������'��k�ʌ�D�cE�S3�����/E��|��I1���w�-��H|��t��w�{���\-r�A	�h�������EuZ|��KVCqKd��v_٨�<'��]|�ń}��N�G�S����g�}饗���ȟ��2S
3��}HB�X���ĕ�³��z+89��ʜ���0R��o�R6e	�V&��7j��`&�Z�������^ʍ�5T�Į�8�
zU#֎��8ß����QW�\dP�7�ǽ�����k�	�@W¬C��
�xk NGGױ�rh�����og=(Q�zWk�ԇ�� &Übu�Rt�'�1d��s���fF��M�2����aÆTm25/�10�W^)0��4=��x@N%אH\SPo͚5P���S_�7-M�)���_���vy*sdV	 ]C�d��ZQ����w���r��e0����6�N���,��,����蠿�7�Y�_b\�ɂ4o�+�3����~Ha��u�]x��<� ��/_~���KB����Š�x�,v^��0�W_}5u���j�������=V�?�~G�܎�����9�m�b����y{pي*��v��8���HF�A�D�  �U�"(�8��QP�DE���%/QAQ$����{���c��;�w�����L=<�i��]�j�w�Z�J�@t{�4���_�袋T�r�*4�D{��:ٌE��i�� l���;��o�o=�ҭΓ�t��O?g7,���U��%��#��1����H3lt �QQ�������=*��&��y�h������0A�-s>�^���e�n��g�!t��k��F�MFʆC�<�C��kS�Mt�Z�u$Z�yx Nn�8�3,
.�ꫯ�"��\�`��|���_,qdb�ؾ�;�հ�x/�u_=��O{5=���Le7�W��W_���Ƨb�����W���e�����v���N?�ǳu�����E*��ox��o�y����u���5��������*
���RPE�ꪫ.����	�|z��E�,&�Ԗ\σ�+0�N��KcPC��u��Ӕ�1D�^�]1�wم��|��6�p��Xu�9�M�P)o�C����)_�>��5<�
����8��-Q��Oů���JK�%��`�O>y��k��|���{�c��d
I�0+�2��b䡷Ke�v7�|3� �ه	.���9s&4��4xM����ꪫ�+���������JB�At�Ri+�oF	���J�4��!����~�B��EbI�`TPnG�UO�����t"���W��v�,+;�sD>����n�:+O�`8��Ë%� �z뭧n=�F��4i!���ǈ�����7wk�Ҷ �s�9G9`M[
<� ����B-���0 8[��_��j ��3���ur�Q!������/�>�͛�c��\v�p��6{����8�W�枕U-B�j�y晼"ݢ��2�����ŝ6m�9� Ucâ�r�)����lW��J��t�Ip�K,!J��2��A���Ѭ���
p0+��
j'����Ł��Np��XD�:/�۸����I���s5dM��1TėP�y���E�@O�3���%��;��?�3���z�Ɏ�"���/0���^l���s����>���)�h���@ZPo�vнH�g��u���	J�y�>�rҶP���^K�p�X�D�<l������O?]�5{7�	 "�0�lо��?���uT��7��w�qX�%�\2���
Y�t�M�����p8$ơ�U������wD���-�9���C����o��FHݮC#5�ߥ�{�9�(?�����s8�ׂۭ���=s}���dN;�4�L=S����O~�4�B-�D�N> ��{|�7��ˆke.�M �v�m��Z���T8���$��������__i�=��vt)��ލ%�D	L��#�J��r�x>
�����Sw�F�U�ӟ��}c����cݱٺ��������}��?��Yd�%�X�i��\���X��~����z�K����RP����~;
�+_�J�*t��ψ��ؤ���1���
+@�4jC-�$U���n��裏��Rk����|�;.��r+��U��i�}+��!�o��2�]�%���}�	'п�e��?�c�S������'�ͻ���3΀&ӧO�}�٭hR�eNQ��<�H��w�e�	W���L��?~�W���[8E����w���,��W,ق���#�����'Q��z�6٬���nm�"�y�]���]�)ԕ~�+����%=��G|��`����n��\j�g������1�a%_B|ƌ��T�K�\���/�6[�2��rZ���o�+W�Ű	��f8�?��O�Ì|X��x �F��_�	Hew���{�3Z��4Ǌ,���2l���1�����Q�f/C9<�p�!]f�e�;9wd�"���K.a����w]�-�"z��ߍ�^M�K�< ��`Q�-�p$,6F��_���CE��	]# �s�1p��h�3V�z��?���<=�p	n�7��<��c��S�Q�����x}�W\q�M6�D�6T-l��ſ���@�o}�[r�>�>���E� J�n:ϧR�{W\q�Ig���|�6P/��׿�u�B����b�aF���v�a��{_�)�M�#�0듟�d�l��Q��� �S��0�����QG�(���*F<����!}�Z�n.�b>�~죏>��o~ݮ-�"�#�L�`\'���'��[�����n�Aj�\�s������r鶑M1�{�|�D UXw��.��O<�De�8`7r�J�n�i��i<�*	�>V��ܭ�a(Q����6]S@�~0[?vg0?$�h��S,)��ͷ��aST6�������?�9	"��]�S<�����n����y�5w���x>��ì>&�TJ�.}7�Y���z_)Υ� Пy��p����S�aݱw�x*57Q�@�k���U+�!�X����Ӕ�I&.�U�_MO���3���Wc�=�[�H������)�R�x�mH7�p�!�:��x��B���:Awt"�;���r�D,  gC>��
���{�iї,K�NIC.o�
��E���~�	�n<Ed��)���zꙊ ��`@��ۘ������෾��:u�QQyG��	�4YŢ*h����=�TA�����؆�~��s�5W�/C1����tn���+�]�tV{��o|���bK)��_4��;�e-`�lDs@���E`�%� �9z��\���e��Z��
��/~�߼����g���s��nu�	�c��<>��O�I1Bf��ŋ�C.���ATX@. .��仟D����*04��so���W����L�#�
`�V6�qy�4�p�``���XW�����p�@�a�c�m��/?�I�?��TA��A�dw���aN�l2�b���de��c��矿��Q���I	<�쳬��Xd]���2V�l�3����Z�ikڶ�'��w� �����V�} ڂ&ɴiӔ���Z�u���>�pP�j8-D|x��>���)�+�f>T��uGߢ^l�m$z-�1g���tTµӝMi��|�r���U���\��oq�R�e� tf�뮻���$�3X�Tt{ꩧå�^���)c�i�p��g6�l�n>0�:^�E��F4T������X���h�e�U$���'��T�P`�S�.��K��s�9��|��_�g�y�؋�Z���.���W]u�x$�(CR=�.(.��ԧ>e��qLϲ
�A�[n��!�a95ץ��4A@�Zk-���+�z9}_��p�~�#�v����-�����/���x�C�nw�����8��v�fKT>�/2��4��)�@�E�SO=����ٿ{��<0�3����'w� �_���'�DCB��*�F�����|�k_�=>�я�|�B���|� nT�̙3���S˱�d�y4 ̀�Q�i�7ϥ�����>�o�ůW���w��_ܤ6e�o�949��ѓQp�HtwY/a�d�vt�w�GR? ��������k+�����FD	E�@�/m��Q�[�#r�t둸��1D��}�Y`,��R^�4���_���/�0������Riҭ�d��0��O�ӎ;������W)8���0W\q�hS�4�ƀW�
�k��@u�x�-�����j�^{���O穪��ّM��߫��p�a���a�\0n�X�` p��0嘄/NnrF�I �&�l�e�{ȫ����lͺWH�l�R3��<��2ˤ�^���h�@|_<^zɱ�-�n�A�]v�e����S(���_x�貖[S�ګ�&��s�y睷�j+���S��8�{������.�&:����]r�%P��_�20���x���_(�SN9�g?�L�₷4�{�Yg�-���6ڈY����y=��C�0���5�!�1e]�B/o���K.��t��g�g�R��#s��j����p����]w��_ސH,�`�ϰ�����?����O�7B�p1�0��%�.v�)F-�y��h���/
��Bҭ
c�s��߸l������#�8t�l����CB� �v�m�mS�Vl�~x4��gh�2ow��dR�ip�`3l\q \=��%��J��-�G+"���k�񶷽�.���E<餓���t�MJ�n1]Pi�=�X2
�[�9<���{᷵h�0�3e�'z�αsJ
�_!#�&Ǹਣ�tV�%_얏lh0�(:����.���ڵ�f�#=�$��~W+BW��n�[L�]�	�J�[h�,�G���-5���/��v�n�5��낭:π�;��s�OK6N
g~�������;�s�dV�ݎI��H=\曒U���o����z�v�m�˝|�=`�-tκ��k�s��y���o}���Ї>�	-IEvh�n���a�kX�1�Ư~�+�2��i�]"�7~�+��x��p�(Ӓ�$���hr�!8<�,+��E�R�?����p:��b�d�YS� ,Hf饗����oKC����z�$���ĦAG�&�<?0Sٻ���0�{<���ػ�_~��ؙı"���P�����|��BHQ/x\M�8h��弰G`n�f�M7�#�7y{�<�����:�[o�U�`���EՐ8�̆���o���ػ"�*�^.k�z�ە��NiK�G(	�����٪�	)�Z,��F9�`��8nCn�k9���@�$V�z�W7�|�-��;�#��(0����ޖm�#s\J~<�s���>���|�#�q�$��aޘ?l�!�ڴ̨�h ��]�i��0?ڸH9��G���v�m�W�/��~R;U���Ot�,����*�,-����-��vԢ�h�����@��σ>M�9|_�S����Z�IYU�BI1�]w�u�UV��y睗� �p'�O�I*��&��KU�� �a�8ͳ�>�v�R�������
x4���7��ю�GI͘1���[,��b��2�����pʲ���y/�3	4�zPU�ysnz$o���_%#a����e]o��XVDIl��E�c�1�^>(�2�2Ր$�m��U;�\s��-o)�&�d�D�Y�.��ՑM�ql��ÏmF��z�$�a�O<%Q�Y�Ȝ+��0`9z�>}: ����N�y�`�T�����9�K,������YP���k��R*-�~@H����c����n��v�9]a�6�C7tf즛n�&,���X.t���^�H����_}\|9�"�[���C�q��<�L�}O-M�=�V$z�����cP�>����2��?��Po��¨
.2H��Ó�Gn��Cxp;2�t��܂
+���X��*G蠃bػ���+��=R�B����$A�����}�/��&��#J=����O)CR�o|E�\�Ǟ^S���;�a��J� j�1�{ad�zW����W�k-��2y��3�R.���b��*p0$vT����^���Ճi�g�}�v� PD��Wg�Q��Z`��!�25�U��T'��'�U�G�����6h��`ŕ���}N�E�	ƈD�
���#�@ޥ����%��b8]��7�ᦪ�&��@8p�
C����?��W��d��ىP�s)�"���ꫯFՠǐ#�F��B:H�,D��p�t�B�S=���&� ����2#de���;ϕ$:��Ж� O:�$d|�m����$�3s�9'c�U�\��<<�؜A���'��eb�X���+�5���9��c1�M˅k�VY2������/�C�Dm���`L1hNGɛv�Լ�#��JĮ���)4��Ac)~p;��U�5�ٻ�J�+^K�?��Y8��N��!mH��? �, ��6Q1T	0�F���޸��P�B����9昃�48BB�ȕ0��f������{0�,�|����\9�Bq;|�r��v�%]��2Z�����0T048�S4N�WK�mY��Uŉ����"���
q�1�f��]
7t���̗UY��k/H���j�G uq�n���5Vc��F۠��%�*�G{����-��B;�)�y�i��@��koR�;�t�IxV-͒@<�(k�,t��?��Ӻ�(Mt�L-��~u�\�2\�;�EYd�y�I����"~��i�9�"�smf^����B[���ӵ���ed�#�c��rXGX�GT��M\Y\�J�,��˗�jՠ��]<��?3�Iٞ���#C#����F:��~����n�a!5l�W��٥�ķ
B�`����D���{�Cu�?��K�ސPS����@�dx0���UY7'��p���Y>;x�Y����aH(ϋ�Q�=hO��552(r���}�P<��!���d�7��TL
J�ݻS>�=Ƙ���@-I�JAN�g�
���R�: �X�����ϲ:F�Z�����˔*{�@�	�`OQ�,+�ΰy�g�b��Z8��u�����/�����|l��K;GQ�]aJ����*h6���/��B:k��%��w�{1���
�dHJ�g)���3l��8pV.� �|�_���N���A�v���E��!��.E�s.4�&2�)�}kxt~��I!� -��t�n�_�im��o����h�A�E|O�}� ��F򠺹��p�V5�|�H����ԝ�=�r��sY�27uU�ce80 6���:�(t;+Y�����a�vՊ�KK���*�I[d�v��B�Nlɂ�ݏ�.�)�+e�Ү�{��E��s�[h���I'}l�_|(*��^E���3��W@
a��VMy��+vт:��ש�Wz�,�cl�*���S���;UE?�TH�%�7�/߶�hwO�ibb��Ѵ�޾�(��������,ۧ�洖��'�9}��>LS1�N�G���N�3�o�����n�S�����O��uhJu?�&�v���xi���X�ė K`�,h�:څ�����`��2l��=e�Lg�i�ؼc�胆�|�z�!�Dd��s~�!�-,.�G�_��)�+� �%B��]H��ʢGR�%s�~�e��Z���2K�������5,k��H�u٤LH���E�.-NAݧp¡���5�=_)��"G�n�6���U�W#�t"�j�_rd�"�Sן�1�r:*��G�L̦�;�G��� 
)s��&��eih�ֿ�H4D遪�h��]� �T�I���s�_�E4�q�?�撩M���Q��Z�N>���Z[�8V��!1������0e���2�$�Rn��L��e�A��HY;G��g���sy(3�ߪ���8�8����5�ªCvM�j��������;�N����O����b8�9���ga����V{�D �?���>_�r����ܰ��|���\�WFyVuy�*d��n��."��c�CJRۇ�(��#�Bӌ��eXM��V�x�܊��QVn�!EM��x���ӳ�
��"E7��<��]�j'��*����ޔw}-PiQQ�����m��y!��pQ��U�0}��)�[?�E��Ӧ�Ťe���nٹ�-M�!�WU�;U-,�4�cy��B���g�\06��|�_/��TŸbD�r#E��m E�O>HaS��}҆��|��e�k<^�6O�Qk�-{�z�5��F�<W#*�N�	����]�K�՚�B
�\>�����D�.��D���y�Gp�(H��g_�+O�֚�z�S��GG�v��HS4��� e> �,ޘnĖ2������x?*����l�'͓��Z8�gg5���d��P��WxA81?�囡y@,-��_�B
It'��O[K�sҭ-Mʠ�E����v�!{
r�`���-T-���g�9�G�| ��a��/�͎\�y�g�*r���C�Z��F��~-}���-B����V��Q�jH���+^*'��$����P}gs���K�\n��2����m$F]�D
?lp#�k�W�N���mB��3�-�(s�zN�����b����:h����o�!x���b#I�$��5aʱ�� Fb$-�����-�T��
��d8�C�*�S��i��-D)��3KmvrY9��^�e���0��o�N�-�ƚ��"0��R0�o/�6�16ji�"j�i��:vf�oEjc�Yj�+���R�$6Cc���v}b圲3,��:\R � ���B�0Θr����%��ۗ��>&i:zW{�tH/g�zRc�j3��x^`L����_3��	L��#�VE�{5�2�ZET�i=֣%/r��w�G��c���A����g�28�g8�BtsV%?lQU�m�7�b֋zy�X��m�o�[�j-\h�:���4⌰&:��b�F�!���P�=��`m����u< ۉ�tR���U�%`c]�(��oL�[����\�{q�
�$��;,#�M㯑��@���e�E��l���;��5c������]�:�Aj<�Q��˅P]��=�\h�㹈�W<�^z��b���@�KDe�	�yuC���Q(��m�f���ɵP4M[A#�Z+����|YU����0��ӹ�y�.�`/ˣ�,�;9��"�7���В>8���32fm��̮�u�����`&dSWB!��8Y}���*�-g��k�Ĺ~(��[%{)h�	�9���(�ݱFN�9+U�\�iQ�Ԛ�Ѷԋ�%���&OQ����a��~S���!ƹ��6uBVBS3���������Ǩ�z�Ŗ)��!.�%�芰��-ޑ	��g�y�7�kg�k?���N"gɮN/礍��>1�Q��Q?��Z�~>%o�ݞN�iQ��a~��a�)����_{M�iJ7ʃ5��]����n�ߞs'o{��Hs��QӖ���줪����c?��s3����7@ո\��t����S
׬ĵ�)0�1��b��T�^�^��<�i���h �f[�+��L���r�}��J!k��1r[��VJ����Y<#���c�#�J��B#%�D�����7v�`<_dnԤkԐ^+�OC�^R֧�PM9�:�ٵ�H1NCn1#v2*�3�a��v��"Y�*l��)�d�S ��v�ͽ��(s0F\�sx�<mGo�{�G���������5�4���j!Ie'$o�:��NL�<;/w�W/�)\���K��oM�˗]�O�>��5�2�uq�ް�D�'-gmM͕U�7�G�oO{l𖃲�z�r��k!2����ޑm��U�Z G=Sذ�+n�&����z:1v�w�����oGRkS'��)�H�?S [�|V'�2��E���0.:~�%�Sf�(�-��1�m�m�E�󙟦�m��s��hX�~��?ذ��V&���;QF:9=R����Q�:�W�@�/-�Ư����h�~.,&����Q�0���nB}e�j�QW�"ʑ�Q� ͟6y6LE8�`����8�K�B��"��{�9sH���5a�H:F�M�ᱍ�\�N(�Rk�����#p2����еW��R�zK5.FrR���ۍe��VM9�a����&�9v�^�0����*�^�
lG�5��!��<�8�ݦ��xx���>I�h�s~� ����>������6l��p�&NHȱr�#�}6X�����GUX�P���7��M��^�ZWe���p�/;�}��{��@�4�Ph֔@+�[��ɸ�vQ�kעF"��P�jR_�ux��{kA�Ԭj����ț0~�BW�v#��jI�^��ýMF;e?ƴ���m�L�Qm��]~cVI����"��75�hi1(��ĉ�ѦNj+n0ƀj�d`mbSV��M
:�fUgM�B�n����Mc3_���]tTRNq�+XV�D�;�ooh!�ab����֊2�;��vBQ?�����i�[j�i4�z��	��ȗ�1`���j�h�I7g�9w:�7���^������́6v���aM&��Mo�������2�P�E'�$ev��9�9�Fq���=�M;�8�C���)b ��<�BPW�����r��%e-�u��P9�u�laAk��|TX���P��6]q�u��Ff���b,_U�>�h!4T�ps4���B��Mͭ�����d4��f�����e��f]����uT#:�Q�X啭��J*���i@��U'�]���-g?�;�3����&ߜ�0�X-D~ń&���Y%�z�!��AV�x����)\s���=����˿�dNK�淈j�x6q�D-Ƽ��{��6r���Gqvi(R�����V�]6�2�j�w�j�!�Ȧ����X�H�³�זWH�EV�6.�Y��r���Gth���[^V�Q(^S��?��-C����J��8NQf��H=�V1��Ѳ��|$��>۰�t6W|$QK��Rr��1"n3WNY���'�R�}�2��0���5M��!t�:A�	yS�u�e�-�\����n��9��Izq�����,�!r㫑Q��v?�Z�����nm�h[�	%�B�1�~��a4<��D#�P|�f�7Ѷv�Y��|T&�+�e��4����=�:�g:���#�┣�|��EG�Y���C�Z��.E��z�W�J��1w"���J$��{�1�C��Ci��i���%��͍|E/���3��0���	W�g2egj�aϡ���?+�/F�e&�R�����脍�"ŋ��	Ix��jr��	K���ϡ��zA}S��a�TӪ�H�iY�ZX+:E޶J�6��E�nj8ˮ�)��!��Ob��jE�G��aHi�8A;ު1[$ND�6uE��7�¾A�W�#1Җ��xu���Q�N{HAA[��-�ǵ[Z/�^�8������	%�:�
�G`��j
G��������b0�嫽��ı��-N�/2�5`JY�^k��,���yq=ٖ%�=X�#�׿�"�&k�<�<i��e�t~f,g4}�������ٛ�sPïfNg5��E'�E��8i0�g<�p)C�<��f�-���b��Ȗ�r�KIG�'���EHJac�U�I�c�r��&E�PB�0wSӯ����ځ)'������ʰM䕵��ð�՘!:�~�潷����7'*��_m ^;�V����V��bhG��O���@����Hs��(����1V��0�Ⱥ!���
����0��_d�O�xhܣpo�����c��O�{o1�����c3��m��KX�p�8�(j��݆�V�������o�x$�O����U�ݷH=��E�6ҎDʁ4R�'6��#��Tu}�:(�1�2�@��@�${N!�����	�PM��O
��a8������M���}\�o�RC�.6���]��v�aV� d�X����b��O?V��h0"8��V&F
�����v����T���bQ?��FR-A7T�d���1�}2�����1�������6~W�t��~2�(BrH
�� �3�S1�=�lw#���4d8����H��H�2Da��~*MXd�Ws�ʰ�Z*�4��ғ-t0+e��Tj/�%pa��Wa�F�o�ٙ\�zmH$�A*�t�!�w���߈��'�G��Ĺ��[�o�F��b���<�4$���"�5;Y��9��;<F�ڻ�E���~xL�'���\5[E�賦���"�2W�|�>E\���;�c5��Wt2/�������o�6b,�z́i�D��tٔp�v
6�"�);���o���
�S��6������ƙ��!���`\xd�8Ұ?t��])�w��$�eT�O��"�δ�	}j}F�4��ԝ����x.����ܕ"�6+sK�ڊ\v�f���0����+���ӭy��CN�x�)lZ�!�����MH�����Z�"2y�x���2K�-��e�LW����*w�ȧ;Z��U�E��y,�@�
|6|W�EH��b�9�{Y�G����j
�F�(�҄*i�rQ?GF�՞$�/B�Z
ʨ+2"�׊kS���y�Օ�I9�5>��TS31�9�C���my���O��`Ʀ��kՓvH�~�����B3N��?o�G�A1=`>��q�k{�9eY��ג��������|V;��U����[�q�&�a9��㜟�%ƀ��B�|/_�3����M��W���nr�d�T��-�u⌀x-�S'�E�U���Zg3���h7�"P�l˼c��jՊ��\��Ӥ[�~�D�5M��{��]N�M^
PHޛ����-u�:���v���6%��.����m��Hm-�{�����������a��?�NE�W{�g������g�H�/B�����o~��Ϯ�MeV_z饿��o�b'���n�2���[����V���s�=W�N�a�1D�(?����d�~��]���(wry
�$�	]�+m�����tK:k0Ն��)��P��7�i�9�x�[ߪL������>L6c��?��U�d*LmT�V̀�5u�Ekx/>`��n�N�2���V��a;��Je(Ĥ���PFUeu�y7�e,'
$Ԧc���2��sN�$����/����a(E��A9�ܨǪ����!Q/gY�BRJ�s�����L)3#��2`ߵix�m=7o�%窬�bH���m`�[W��h�B�Nu۝Y�ǜ���"8B�;qk��r�ϖ�2� C��6\��%SS���~x=N��2����¦�|���9�$L�g(���(Əb����W�(�OL�uB��4�:a�H =���ϧ�D�Y�4s�~�]ekTË�gUW�jYUk�q�,GvD59�����u��Z�c���jr�h�%��躌�S�!l�xX�k����}���G��n'��%S� 8YTW�@p�?�S�$6��b}6�Ͱa�Y��X4�v�B��]�}ҥg���-L(����bk�^��!��&�`
�*Glc�h�l'��{?�>�C>��wiN���Z�z��wG6�x�0l��陕��!��蕵�Q
U�4��+G���!K�B��ٿ�Đ��������4�5j���g���"������9�ՎV*pp�x:�4H!����J���!ӻn�ٿ��|՚=�"ߞ�I�,ū�Mݱ)�w�f�c���(
~�n�W��o�{_~��W_}�UW]|��U��w��ݭ��z��7�w�}3gδ�oj��La�����J+���k���
-����+7�x�M7��+ ���x(T<��x.��%��E]����+�L�hC�p���3f̸��k�z�)^ԭ.
��M-����8t�*��A�"�,���Rܕ;��=���0�}	A�&ܙ2�,t��r�A������|�;�7��뮃����'��o'c�deU��e�a�묳�ʰ!-�>�(a�?�0�"n�5�!���KL�6��62�0l�d�7�pï�k�JU��i��E1A` (����>Yq����w!�i��[�n�0v�'r�����Q5�l�0�}���o��9�(fM�U�M�������w�y!ԆU���s��w�_�;LiÔ�y(#9�g�04$��o~}���zVQJ���)������t�4����szx�j�$#��o����3�|��X����&k�����.��.6G��9<������8KmBn��*�����&���s�=Є�d�
ޔa����2���S�Ne)?�������|�G����+�~�!甡?���YJ� JL�7Ї���g|g�kj���^[�A%�S�b����.H�F9����$��];^���{��އB��sd��+����{!W

d��וs1l�1�
�E7B"�K���Q�ٟ�	����.� J�`)`H��a��J@��P��ŖQ�'Qb�K-��MWRÍ�]��*Qj�sܱI��D��Dq�9�X@n�&�$ҊK��v0'��l��l��F�:�ğ���\sr��c�Ap]e3>�,��&����Y|���Gp 5`�E�9�F�&=��N3rf���]Y؆w=�����+���<��+o-���?��p#��*�Y�F���0�I�D<�#��Cհ��J9H�3>�D�B�MQ�!���:�+$Xk��`x�3�\s1�^x�� �$0i��ŵ�`���7��)#g����1x��;�d�b�_ c�Xm�ՠ9V[(�d)�U �e���,���<����0$�Y�^zi�_b��y�h�Ib��D&�}w�R�'T
���`)� �b�h-�r�-7A����c���	�@�#���T�a�������rK"*����0:���N;���;�8(������&�@Bٽ��0���=�z��C��㎗^z�	'��Z�츧f%.�� <}���v�B�C�~/�6�dF~�i��y晬�uJ�wK�Z$^[|�S���G>Boa  e��6I�t�I?���ц
�9��B�$�a#-[n��aG?���^r�%�sdO�����c��;� á�5l�ElX���_�s�����G?B�75~��
���{�'��1C�T������#�����B!�\e����Moz��d�ض"���3�Gm1#t+þ��+{խ�{��^z�җ�����w8��o��v�ٓO>��/|��`�0\��aF�_�,�r�Q_|�'����-E��}�ݷ�f�ω"2{/�0i��?��sO9���5a���Ʌ��{�'+{C�U�G9 J���O?���ћM�C:)�˘`�u�]����$<�g��0u�Q����/G� \&y;�w�Y�M7�TW�0UR��g�y>��!��]v١��F7Yb@���!�{��G?�Q�����c�P/�#4 49�3�nM�1Mp�g>�F�U�.H�'̻`Bȅ����ફ��&�gi��OX>���o,��u�F�1K���z��;�K���l��V��<�[o=�-�K0��,@xp�y�}p0^} >��z뭡 kJմX,
���v��'?A�̜9�5��4\hB��D�l
@�6t�~�<#G(a�ztћ��*�β��  h���1-��}�v�ͳ�۲�G}4�]����v�]�Z���U��)�?AmL�����K�?����e�]P��D�*Fb!x  wjմ7���\m�C:��Q)��Z���?�O�~�ʍ��p�K��%���a��ZT�Ff��b�-XYd�a�Ɔ. �5�,Q��-J`��IYL��6@�@2���<��7AF�W�Ռ�@��Zt��±�*�z�E~�᯼�
n�$�[�L�1@
�{ǆ��\rI&�S��9�$��FW0�F�0ʼ[^TI�v4�i2�P��[��b��	0��N�T�������h0u��-�^L�!@A�#�Ƚ|���¨�������n�݊�B�2`X��	�l���'ft��y䑿��R_Ip,?�jgO߿��ߊ@������6����@yH6��� |����v���+�刚�3G�t�A4ei�������xȽ���� F��HYe��[��7������PJ4k�L��8_��ӝp�id�؂�P�{,�Jy�V��r��;���|�[ߊ�w�{r���<%��җ9�DL�B`�����GI� �wE;��7R��w�@s������A�P��~��Z� ���E%����Ȃ�8�S��аM�� Ԁ,�r���?�ʄ��+�4$��#�����v��|H�����jX-�ǅ�qha y��T�|Vu9���xKӂ�b�L�ԟM�PF_��WQL��)T��B�۱�п��4��p���(�3�B1�������!K��i�%Q�B88ѫr|W^yef
M$�e8y"����k�	MP^P�1I���h�U�%pD����M�� ����c�z��aU����C��� Z��pO� 	fo�]w�&h ,�s��+�<x��7�1Y �j��4O��%���u������7�{�N.|n�F���j�P�t�F��+��\^>��6� Ņ�y����q����;�X� �� R�l����9s�̿����`����d�1q�,�dV�t�3�v�Q�N�_"�DX�x��ӧO�����	�5!�W���#<�n7��#�[[��w��]4�"�8�0Ȼ��M�F��$���tF�M'W8��H��N�����������O�S���f��1vtn�����|΢�|�A�KK4��Z�B�v����"��Ҽ�j,�48�Vݞ`��=kL�� W�7����D"p ���`�O?i��1q���F�>o����"��w\�-B�B�o��f�1�e'��MU�c�x�*o��V��;T�ox�_N�y�傪L���+.�z����sW�p��O(��J+�L��Տ,�V��+��"h�������H�_'�g�,�Ґ����=x���o�}l\z�:Y�C�8)��bՔz�&y�n��?�yV�͘1�+R�E�EVb���F�p<�:{&D��A���#W;~)��}�{߃��ZQ�  �k����������f�����*�TN)�A��:�N>�"�M�T8Р/�+�.B��5�A��{���_��r�e>*�Yw�a�2`x$-17�Bh���W_�B�[�)�ϐ ���V[�ZO2�Ֆ=�O#3��Z��5Yu���JvdC���N<v衇�$��f܆��)�7�D�8�NaO�f և��5|��/~!��<
Ϸ�x�04�R�[7R(±?>���p�̽��+��L����_�����[r���5<��o{��D���K/�4����	< ���w��+R���҇�	�u�o���hJ���_�>�H�EG�w��ӥ��"��U����?>���hz�R�����}WV����y唫@�{ �l�}����F�TܢCr !��:�1��\�7ܐ�w��]���y�t��!; t�u|�4��1�J���p������NN")�j�&U���ȴ���?�۷�n;�QD�����*H4�B�H��y�w�%�P�^�O�()r�zD�+Ѣ��lx>��Cp�_
l��/��a}4'Z����~&{)��kI��c�1^����G��^��0�<��ӵo���di��5�b"��W��b�-��CL�6��뮓�Ĝ���+du�a�O9O2�D�[x#h����3g��^M-���O�kRP�b�$2�W��=�}�CT�ǎD
�ai~���o�M|ة2������|s�Yg�G��W���Bf��Y�	��o��6�|M���,��QG��:�ȡm�6U�.��?��|���"V��{�����bE��c�{�1��D˖����"
���ƣk|�z$�Cɜ|��
�5��1�馛b.�'S�0���x/���;/e�j��<%z�S���4� AI�]w]����3�(nh�I��'�܎�ȸ�s�vt �bRN��������ٝ��m���c>z�欬�����L$���|���<�W.��|�_��'>�T��?�e
,"�0��<�Fً^>���o�*4dA�ˡ�2����:�l��:��0����X!�9�'܎�{��9�Ä�-|>�R�v����K���H!��O��m0��E�E�|�~��qV@"�w���@�l�����mL�q��U�I�������7Y��|�2+��#� �rZ������x��H{6��A)�y�^x��o퇸���;z��W���A)�����p�A���]2�H8�^�(���=�������_{�w�yg���/��W�u��j�>��Oo��&���W��=�I�G*|}h�a+B�$�}��r���&��^�b0�*���.VK����s�=M�^�['�v�d*42�ɘ���ao�����"�Wp�����Z��4���eH��	f�J�[�D!��wzvV(�n��+��4�.�0<ӈ�50e<�裀]���)��hY�=$z�6�&m�ۋ��B�	w�u��_����+�Zj)�&��\�)邕�n��0tL���|�S��;Bp�lL<�h�G��SO1�_|�0C��e���U�X�J����jt������g�y����m��\x��m�{g�~KQ�[��  $���G	LɗY���1e~��k�ܑ�U��b0�K����~~�%�@4 �Zk�G<E+GRvl�5�Pl��K/��D��9��B�p<*��=�	ׂ����kɨ�cƚ�%���z���b'����3
+��3f���/�,b���;5v�i'Y�&>OY��� J(����7M[!��!�;��2JG������{�WZF"��4�r��Iko�/`_��7�t�i���2 ��>��E]�O�:ո���S��Ӱ�H��w�Y�� Qm�r�:ƻ�<��5�\3MԴ��,����ꪫZB�ڽ���~�>}3��N�QIs��Yd��|�3�\s����);�Ƽн(=��a��Jr��6��q�P3K�g}e���袗U�rv)s��{��v�$	���x���"�x@�9T�2*p��{����t����>���Ƹƃ���}NW��s�>(	6U��,Ю��n�K�M�~��ϋ҈dj�֯�T�x��[o=��ǚ+7�{  ��~|҃�ТH�f\(�������n�_��j�i�)N�qbg+2��P����+�/��g���������Ce0�B\��9S'ܯPS�Óu�NE�����x��h��������?�|򓟼��U�%ҹ��E!cf����{q[z�#c&[�Z~�Ὢ���e�7��r�4Lx��]u��z䝜�9r����կ.��2sd��r���[���PT����QI�r��O<��
����b�uGʣ����PL�;�|���`�T���L�r�k��VL���c��t{��?/b�ȇ��zSLN9-���[
�-��6{�̐�e0��g�;�䜴)��=�1(����H���_~��7��A4̂0$d���U����:w����0�>x���O�:�v��V�jz衈R�Ӛ��!A�Af�d�d������Wz���)T'{���'��������$kJ.�	�`�n���DV���>���$���R6�6l��
��jj�J�|zu�^��G?
�pU��/��@�{�'~f9T��P>U�r >�r���r����ÄͶ�r��?^@4G6R�C��C�O�=�ڟ�k�!C���M�~.m�'!>cK��ޖ��ʪ �A�����ٯP�S)����܌��f�' �9�C�O(M*�t��H�G^c ���Ѿ袋P�-�"����*H�Ϊ90Ѵ����/`�+����s�#�;5���:L�֜̓���� Q'
Z���#�v�my������]���Wx�rG��G�3P�2u�b���%�v��c�1(�9l����ToG�ă�
M�z饗��L����=c�b�-�����-�t�>��]`�0��	v`v+���7�S�w)����� ,��ɂd^x�8T�b�����`q�%�}0�2Q/H���oJ!��CtA�ֱ�Q﷿��ػ뮻Gq�)'σ.V_}uY
=��i*�A1<.!����n���GƇ�g( ��َ���Rlǈ!1pĄ�ȝ,��b�Bk�m����:w�j�J��ҿ�.�p#[NY�1�@�{�G��#�Ge�T,�ݺ�\LȂi��� <���Emغ9i۳��fYe�� xmX��;!��N�
�I�y'ڛn�����-�s��Dԝ��	���7D��N8"�1�`�;2���O��V��-�,
&��h�@�b0�7�pÓO>��xe��ԶFJ:T��7��<kCv�^ӦMÃ}�G"���T�<�w1��P������������O!#Y=H�0k�s��DS��ab����+�������|����#1I�nc�zo�1z���dQ��}:��.DE�G�1����N���o�(�b=��)Buip�zdӮ�&�8���\S�ъ�,�����*�H��⪃��믿��������!��#���p�]5ˎ>�{睫� �	�|�}�Ֆ��a�佤���*(��6x�;������h$>�()3A5�� L���1t�n����J�����E�3Ƌg}cq�۱Jp��}+���;9�����j��E�"
�a���馛n��e�ܫ�c�۵^-DVƦ�j�"��sΑzn�{�_'��w�4�ĩV����'����!��bOS^_4�}�qǍ�
E�u;8r���Jf0�����
-�r3f̐�&j�����1�&ܟ���E�)Tk�q޾��C">(C�}$���������(��� t���*{֛�-�K��zm��f:*fmS#�|Q�t4}J�������i{*1�t�)[:�)� @ED<��`�xʷFȻP�Hx����!<����A��[n�UW�v�I�1L��
�v�
Z(I�L���M!n���5�Gg�v��O<�tLTٰ��G�P��=���:R+��� ��T�s�D48`�yѾ9c��7�T�o�B��7D�RPXft%����aːD�����ݭA��$��NA
�ou�e���0���A�a?��O0c����˗��!�*i\z�Zh�2�mc(2��R�s�9�.�O9���°S�8T%�����޸{��s��j����!��[cs,���
b�_�B^}��N8-�� t��1��x�/M�	d��H�C�:�7�Sǋ���FeN���I�B���^�1�ݞ�:���d��|#��T�H�K+,�*G��D���	��+"q5�Z�I?䠧l��Yf���W^IYB�
�����#�>8�(%�2JqA��v�mq;;Z5�!�Vu �v��i���VgC�Zj��3gƿF�����/��5:O��ky���\�^[}�[���fˢʕ����N·������<�L_6��3����8Ǹ�瞡	l���i7}��曏w���md��ޘb������=m8�{
|����,�]���\ ;~��B7�u�%���uB"�(��ڣZ��`�D����_K���j�p�����JRDme\P�l��]wݥ�N���BP��2�Dj�i�Y�Qk�)<�Zde�clb�ZZFQ�	ils�=7�K��ɠO�FB�u�Y��O.�ɍ�W��T��˂��*�l��+�������r�����yt����=��� ЇEu�p����v���Ձ�E��#7�yo;� v���3��Bf��R�u�L���퐴����7t�/�H��%8~��b6��q��h��Z�(�?J��"���sԋqH�M��{ȝꜴ�X�0�2uݛ���K�#�V3�v/S.�ީ�8����}��E>�_�8^���l�S�K�h�9�:�,���x�+�v+�����e.G�m+r��U�a����4ʲ���=�C�8ڰ����������bJŪ�2�*�-��w��eC���.����%Q�����l�
�x�;46IZ�(��b���U�(���6�R���Z6�T�J'ܤS럑�vU�w�/�S�5�`̡�,�w��,{�B�n>?ğ�Y�OX �����Z0x��%0)�M�盕0N*��9qO����3=c���~���
O�$�V��+�ݢ�:U!TD=D]G�ڛ^ʲ2��Sc��4S,"}`�(�N8��O
z�?j�ĕ2�(��%<e�!�g�y��
����@�X]%q;�ti�L��nu}=�pJ��Q�����Nb�}�mí���ɅF�ak	�^�O���b����t�=5߂���N�qܹ�����$���v���?: wϔ��"�Q�pU��ڊ�Rt<�������H�N.��[@��H�N>?�t�)F�����P i�|�6�_��!��/��z�S�N�a-�W��c՝!v�������;O��*�ad�I0��7H��G�/�\�I
n�s��d���������O�1�r8��1�F�_ij-�Jm<߆.��TrTSM=�	�������!í�+
H/��(X�#6�y\J:��t��aM|b{���?��Ԉ�*�(�ޯ��,��|����Uf,.��$����Y�Nނ.�ӄ��p�<aHċtZ`���1�<#y��mɺ4�H���&>I�,=�Jd�Z��RN�K@]@9�i�9����j2m>r6��W�B��v�W�m�0�#��
��]WRb�|`��iiz��W�$;�0t?�Yv�M(I��lq�%A�2<U��h�d��^��X�:�M�Ȼ�
I�6<\��&+B�+p�oS����� �7�PA�u��eN�ʣ|Ķ��f��<J��p�v�"��E�"DHP((qA[��3�iȭ��6�
'���;����*�����3�d�0�
�֚��&��Jj� �ەp���
A���"r�
��}�h\c�Y7>�/�<z�d7�_خ%�g��j�\
\�\R������9�&,h��G���ԁ��(yJU���{�� z�7OZO�M��焥�����jM&J*��GZSuԻS]�-�q��-��4)J�g�����s:wLNߛ�]aC$�ёY��*:�$"s��<��ml�����ϴx�U,����SL.��qZ�{=�2�Tj�u	�K/�T���/����k�\MH�dǰ��j&S+¼IS�(�E���a
��C;r[�f�$H��\�\�� E����&2i�>Q�;IJw����N�ur�;z�>��L�j���暋����=�S���#�޸sZN/�(���~������4� R�as}�^>�TV�J�/�B�K
�Qz������%o,�s�I�83�{,1�<
��	�6�N� Td1Lqi�s��HV$"��`v�����_�È�nd�G4֚��w�J(0�q>��S�PY,��F+[��1�]/Y�2oq���?������Ԯjl´��:��^��Ⱥ�7�~�a�J���Ć��^t��FM7?�!e�Zp��C���u$wk�
����E;p&�͵V���VD��Ԭ���{��ڋ��o_�۲S�x����kh�NI��K�Q7EK�C6���^��FAa�^�γ�H��Ђ�[��+H�KyӐ�^Vg�t+k�+�ʱ����~����W<��� O��	-Ѵ[��j&��"_?g���/)��e..Sע��Ԕ��T��0K�zj@��Y���j�� K�X�=�Zs	��� ���q*�4f�ƞ�*���kԿ~]�*C�a���0���n��e�@ڪ�p<�"g5���8�\ ��e'��w��4t3�N�ȯz��T�x�'y�)h��`�h|ކ��C�qJL
Gj��˼��CSpZ⨊*1C���-�Gi0�{5ޖ)r^�����e����|9�/�x���Z�ny��WA��P3�6�?��]t��pT^M�Ի4���O��-�ӰP�&���+X�7��MP	��z�,c�d����o�@,���ڀ�JRs�VE��"b����D�U��sQQ)�"�<.���Z\AR�y-��9qX׾Md+�����Lo\��8�E�>������Ӊ��43X'[-���`tՑ�h�7��KUE��1K�<�z:�:Fp�!U)��=-�ٽEa�O�I�S{�:����R�U��/iϧ�@c bd��+P��d��N���TWd
��D�)��S�:�pBw�"���+���M�4�r��ό��o-���S�`�<��,1��^�q�P�7���zJ�p�e�:�i �6#i��r0��K%q�\5�[H��q�\�2���s�[�&&�|i	Zz,���:'&��\�iV.� a�����Cjn���N��IN#���+��b0|��H��	�/����0�r�Qd�"�h�(����x�N8Υ�;��5�z�gT�{�D��b90�	�k%��81r�L�Z��B\�"?��_���?MɵSb�����/�*P���DǞ�Y��SO=��˰٭��>�,#��~���I���\�6�#���l���hE�C�Kx��>���"�˗^zI�HC>0)V�trI>?V����ڭ�(z���:��'S{��t���He{:a�]�W�k�"����?�1@`"�M��*��� #���&,ӟ����3!��U�B�R$o�=ӵ�M�PzV�(��ǔ=f��Ѧ2��GR�K���V��2d�����;+W&I١���3O���3g��1^;�y	���/�X�8�&���.��0�Л���sd�ʔ%��V��4xB&2��>��ǉ���j)k�|��>��z��_#{�vީO�/*��"�G� tn�Uw�.�D���<���sp=q&z��Gc��ri|�G$�~�c�Dh)m��`���~�iq�xU!���<����-��En/�u
���Xt�E�����uH�	9N#�_��K������ٶۋ~Nl�V���t��8�V	�ּ�-T�:9�5��~�Ut�F�� #�*�����F�'�+�՘Rc�~ut�2���p�6ESk���,�	]��6��C|^�-�c���vA�C��w����������Iyo���H9�α�<F.ʜ+�_�d��5��wa�'�m@̯���։.��ѴL1�:�+v��f~��6�8S�*< ����쇣>�`&����#@m�{J����\����94�-AX}8ʍ1��Yz��b���us
}��;Gݍ�����^9�����]�n΅�3��r�� ��7��O+�"�g����t��M�勁k�1G�6b���K� �B1!E�[L`''B���ͰS�9XX���L��X��T��tO,�\Vkܼ����[�����m����o��^�_�¾��衇6�d�~������B+8�����jK�4�Tr��%�����j�>*��7m13/������NN�Ig�G��W]wu�m������FW"���k�XK?�'��۴@��-��R��I��YVVc<�m���!��S�PK�����'�_�g�Z
Q(�N�6���rì�o|~@{>|~�ǔ�h'֫,����q_�ֹ�ס����k�mQ��%����F�adS��Fi#�����n�馝�pD-�:���%sDHu�θ֢**!<��K�஘D�>+�n���'� �u�%�d�nҘ�E���L GXʼG�
	��0e3s����jp�G�[��j�ۿ�ڕYh���!!�}���xt���[�E�BXԨ�S���u�(����@k���X]C
�_��9��u��m�wE�����-���Ң�8i��@����6S��;��/g:��SO��*yT;H�c��*ׂ�њ���19cLM���.���T=+����|��X[���|����s]T&�QN?�)p�t��D.�#=Y[}������pZ��|91$z#�����.c���A��z�#�RR�6����~�� F��bt�_���|���V���<}���]DSIa"�r�Ӡ<zl�T4����ur��~(����oHC�1����!��"H7W����p�&��rj�Q�p?O�f���b�2>��SbRXR�)]�<1���y�{��	]�)���K; TT0cd�P� ���e�ٹ�\����7Qz������	�g���V<�����.�u�A�0f.�B�x��@e(r�UW����[<#��AĖ�3`��>�1��x�1�F�뮻R�GˡM�yK-��&"��������T��}vB1�@g���ʽ���B��4L�:�?���k���{qt�3����9=�|�nH)v|�t���Qi(��35E��u�Ջ/��wծ��J�z��A��Ű�7�|�(M���'�r�|t��Hԋ�?���w�y��P\>c��0��*|�7� q��X���g�]l�Ŧ�������KIb�g�Ug({'b�믿~��S�`���"_��Z��{���k|.E�e�UVY����M�䘨p?4�����0�1�w�}�ꫯ�2��ȩ�.�deuD?��Z.����ov�3�<[��(D��;T�]&��,
î9Z�|~�F��kq���9�#|qY�?hN�����~K��<K�D���K=�YH$=�hn�!���#&h����D���ƻ������)��
�*0k���"�ܽ�+��v[%�(WD�!.�uZ�D�soפ�H��A�Ya�4`���^
i�F��dF���|���&4a�@��٭6��􉱓n�I�_A�0䗾���O�M�w��q�ب���XGh��:��V�mS¿�w^�C��'��h�3f 0�*�)U�O��	F�2�[�??G�bXWZi%o�5Ǧ_1��X����.+�(��~���������:c"�$��b)I����p]�������~=�eG�9-� $c��K{�l�ѫ�\r�7O�C��2o\ Ű�z뭧��\� ��= ~��ʜ�4+Wp*��:�l	���4��g:"&�&��DG���FٗkYJJ�g�Ф%w���5�\��V[	�4%��~կ�*`�"t��nпRQ
^x�?�a9�Sr�:?l.I��1����,���vꩧx��� �H�bS�_Y�SN9E�#� ́�`�Ru�GK��~���g���_~�������{m����T�q��J�`� !�O&�z�3C���g?���P�����_�:n+�W�V�"���Ƌ���b=k�b��ޘ��DA���D��������+��w�ٱ�D+�,/zc�#���`Z��k8��D�2\�ˇ��:��Oj�'>㑟���Їt\R�v�BM���
s�'�/�п���
1��ﾻҸUD���>���_m��~��5��}� ��l3���$D���2����C�~�>���h�ӟ�t����$�#�����C����,{L��2��R�0��O:餖�-s�	��+��G��c~�ha�E.U�2��oοhō7�X��h��w�ͩ��dl���J�G��U����K/]w�u��gW���Z�O���_�Bi���k���J�@Ko��ε�7��MY�3��/��Q�����SO�q�_�����\�ݲ3�r���`��O>�����o��3	��������`�H����.�"gF��\�\�k��9�҂�͉"/l�Ӻ�|�J��<$&��waL�<�L4�cM�E/��{ӵ�̥�>��e�]��6ی�Vt��4�)J�YM�AH�E�N�jK�.�
�`qH�O㤠�X�_��WӦM�zI��r�ؙ �ngA���k��'�o���ɵ��R��vp;��������'?���56��Ҡ/m��]�q������"�B��D���X���o��袋�\�~����j�UCϋ/�x/��O��9U����;ߌ[�q��ްY_KY�1xaQ������t�{~R�S���r~��,�0���N� �D���5	�FTÇG+.����&�rS
ᆪ5�F5:��0�� �|�odsЄ���#q��_�SjW�o���ݜMQ��V>�u��7#	�ekkV(�����z�ᰟ�:�b^w�u-Ö��~�񫮺�΃מ��^e�����?|�ᇇ�q���(��{����n"#z��;���#�K��d�Q�`h��*'������g��7�L/����h��2˨`LЊ!�2[��N;_�R���0�� -��RK-�:����4�x>���ft��1p��j8-�[#�E�HK�A=�z��7�lK���[`0 �L��]�9�ݛ�0l\�(�/1=@r���2R��%���8O.4c��͊e8�������{���x�y

��	���/��++>��rFQ���ݗB��p ��5j�M��ʢ
��i���� ��T*Q<Wkp�1�C.����&ųӥ��𩧞
���DΌ���￟	��]�c�9���2�wy?P��ϑ�-e/$��v����)�����
�+q���闑�uO<�ĝv�	<��fod�`�F"O��l/�F�MPw}����w*�ݧ"��T	?�i��=�^� ��AK�R���g�f�,n�lL�Us��w{��2�mF~���6{ｷ�<IN��-�և�����֥2NP�;h$�}�M6i	-��T�O�W��Q�� � �>�x[\YAOxF��\K?�����r��j�a�~�ORU_�;��������?�'�7m㤰�nn7��  p���-��ۑ�W��GI��n>u��Y  �(IDAT{:�aˋ���I��MM�X{�35RD�o�����C7g��AEj*���0 ����d'��8���_D����Z��v��f̘q�	'��o{�۴E \����>�����n�`���yݎ��z�S��
jդ��[k~V��}[H/Ts��d�)�e�N�`t�L���&Ŋ�T��l��3x̰:��&�+�����;�-^��
H��i�B569�*�L��ZZh4 ��}�#����rr6�9��#�sN�O;,v
�̖��T��`����J�A
���QGq�|�ͷ�BըV�Ц��
h|���sj�Ht�ϧ�n��&:���?=�����O�O�*1)x����j���:J����b�d!Zbl�̲}�[�Ri�2kmc�L�;�5n�ԩ����7d��Ew}���-5��YS�� m[l�"li�f�`��S!H��'XԻ�<�y�ǘ?��G<5�A+p�"���������q؝*�3:�  �J+���"��\�E��Vz�(��񵸠Xxv�Y�â�.
��M��|rz<_f��+���#�`qY�n� ,���%+�B�,���"���v'ܳ�>�Y��#+:���_��v�!MΛ��U~� �D��aK�0�+:%e����ӧ�-�4��Э�y��"�GK���q��<�����oz���00���r��1Y=��^{)[�F������(e,�j)8�3�fs�[;QK,����z��� AhUw�@|
1?�C�h�W������^�MIl�0�R����&���4��ƽ�ܰ��n�B��z�`�aޅB���A�����k��5b���3�@�0�N�~�B�$s#:�����)o�(�� �x���EVVZe��ҕ�쮤j+��K.�ە��}
:*e%ɰ�	ܮ��~�f��"�;�����+����[�C]��1e̬l��t��e�p���$Ge�?����~�W��EY�UAkO���Yzh��QpD�hd�"�\��
+��"u/\t8��[�R)�������D�`26�h��\�ʵ���!49��tP0ealGQRe�<�XM�6MY�M�k/����>�cMˡ�9s&J�����H�`�a�~N������k���w���{���oU��S�cSoڧ�k�*��uv����yx�e��r�-�/3'w�[К&4aجl�\�y	��駟�CC��[n9��/�c
FG��;�@����&Rc,߁�Ձ��x9��Cf5� 	-�J���_i�
˔�ؼ�������e��p)�d�-�(e=�n�O�����������{Ϝ�z�w�*(&�,"$g�$((AEP��1�	�k@��b g%KP$J
HP�D��֭z}��~?�����5{f�y��[o�q�9{zw�^�V�^����4�BK��[��[N����X��i^���|�_D������0�����k��կ�}��e�:��h��~�s�9�nVq�5����Om���3���������L�������]��yn�@��nql\�R��w߁��uvf�	��'>��������Wz3q�aSx���&{��$�J�p�A�z�֧�ѻ.%9�lؔ}�����J
�i�t~�y�)��o
3�Y�77��$3�yF��,�袈�s��As�^W F�Q���pI9����͟J��f
����nM\�ATj�2��N���=��h!<�V��o��&ROΏW36eH_�җP3Qp�|�
'�y:�����y�k$�;JjT� @��駛nr`L���\	�z�)�>˄a@4�|��l�[�;ckD���;Ｓ��^�v@1�8��S�ȉMU�x���C��7޸�y�%����	!Ӗ���V���aF~%rj�@p�u�ϒU�.�pV]��o��A��\����܎ܱ��R��Mv+��� ;�cIWp�I�[*&�k_��Q��A��b���Q�/~񋨲��~^�Z�����!��N�t�e�ւ�:�����q�uDx�3�KS�J��F��Ir�~���A�s46�t_򒗈�*�O)�&/؊�@�+2۬^:jUŹF�d��MtY�wA�)�����}�{?���r~��=y�v�ͽ<�^+��[L\+d����n&J��>����EХ��e�M�h-�H!V逶�6� >����whk�%D�_���J���[r����t�/;�Si�}��F�	����k�Q�V�"��۷�j�	Z�ל��
`��:\/��J��l��nؑ�Ű�vRo�0�9R�Oe�g�r��	BF��R����0�1��S��l�[WR|a���x��?����v��/|�@�{}@V�������m���R%�]t<���~v��6���=A�6���X��/�|&n"wjt�6㐟��'�J��Ld��IX�3��d\g���Z�c�p/���y�{��5���&J^�&2�T�
��=}��ؑ��,>x��.�t|�Ʌ�s�E8�e`a���w���sO �x��܌	�Dѣzxr���v(I��]�,�%�\���b��Yg�f�1�DN�?�xxZ	O-G�-+#�5�8���o���[؞�T3� T7�t�Gq�Yg)�=ѩ?������x;Pf�%�P�� ��f���C���[u�{IAw8?]R���_d��~�a�A-����w��<��I'�����{����3���Q��*�9:FCoj�x?c yw�q�p,kդA[{�ì�J#�2ɌK���g�}V[m5��Uq	��o���*��a{�f�ُ#��̻��n� ��W.�ྡྷ���{/���.��Q�Id��Z�0}�/��^zioy@| �	'��,<�*v3�q���x���뭷��Z��fC	�y�i��𘟙t�_��^���'�ux�V�-1?|W;�NF�!h�ZB�j&��;P�7�p���Kb$J�E�[�X� ���)�V��䛧a	8T���,S����ʓ�,�lo�QG6c��*	 e)}�`��v��B�й/���;9T��k~A:>��O������+��r�� ����ap�e�]��+"d�S��+��㮻�ڪ&$&�f����!Z^���zzN��p� ^a��ˊ+��ܛ��5 �i�"��YS�~�\q��{	�Hy�}xoI� ��?.x��W�H$��2Yy�M+��|��F���w�� 9Q�Y*!�(�AO>�dm&%���:ey1�~��W_}��{�I�L4���n1 ���b�∃0�A���],c���>��f���3qմ�Æ��ޣ�>Y.I�M[Gӟ�b�D\]����1�q�g�oqR<G�&�U՜��!��{��^��W�[˰�$eTQ�ٛ�hJa���쇟�O�}�e�-�QY"�O9��?cZb�t~T.ӛ_�����>��sQ�_�1�%�VA@|#/�L
B���F�n�C���yzR��\�D��Q5)��״D�Wn6�?C��6ڈ5�seBFW G'�x��1���F�0\h�+�n׍Z���C{��GYS��u�C�c�R:H�zk����yb(�#z�G���+)DR��h�'y��t;�#_�)ˎA��lm:���60�@U��������1}�+_I�r]\%��c��	+��^�nb|Y�z ��_w�u����ZJ{8�V`���@�H.��E�ya���wd�Ə�я~�����u�(K�@�9��P�L��ʣ����f<!�9���e�*:�Մ�Q��֪w�x��8��χ�Xu�Uцt.�W���ńKU�_�������=��2R��׾���6ml�%Y]l�UW]�X� Uӯ;C�j����!����P�T`	<�%F�DV���-	4Ys�51?�D���)c���w�}�,��X�籵�d���Zw�u�_~y%���9��2?n��Ov�%�����׿���g�_f�eJ�)��>x��_g�W���$��E$�t�5�X�����W\~�����g��:�GG����T-�,p#��.V	�>Tk�-�Թ��VZ	!e}q�2���Lܞ���P��7�C�^z��d��֓Sİ����t��i"x��71�T�+�
�EHWYe��Cb,Q�W\q=K�d���k�'�N�#e$�*�
�@�ܭQ�%6U�m�+����kCm��j����CD	>����4�f���ˁ�@:�&��	K����+���<�{�t������E]���]�?�4U�?����7�S�cz��qX(�s��_	{Z��P���tꉍW3w�.D��A�)e���^q�#�����0n�+^��VE��	ڌy���uۣ2zw=�<`��6<�(1f՞g�����I�W�w�_��޻��1�9x�T~K�$ס9�U0^���i$R9WU��'�ރԛo�9�k�E�sFN�,%�� $���2	7��l �B� m!�K,!�B��-:��C�Ϩ�vT�J�Ta/�vn�&z%��`Yy�Hq|�$9�#B0��]8_�#�,:�pH�ѹ�6���Ձ�a�"�~�P���ک�;X�W�sƣ y��M�uUO�s l�{֥� ;&I+۽5m�H���eY�c@G�s������b��qG��4���s�=��h2/
̓d l_��n?�Pj��)-q�&p#�3f�G����-�62�Ț�u��o�"�Ř�w8�o�1��/
���(J�N �h�f�Ofk����n������eU�k3�u��t� �I�9�I(��R�J����4���ٰ�9���i�Wi)�Fdk��Q�9�j�7ɡ�����ԵM;�cra5��5H�;�1�85�_<���+cA������Z��TX��$�攉���ad��y�i"A�cL
]�/�]>�\�P̑3=iw��&~�����i�T�[ɹ���Zt�QK輦i�qȥؿ�S�*m- ��w�f �'���Fdc����˺�B�A| ���(�0O+5��#����_�<�m�����z��F�q�ci?�6�8w����8q��k���6$�%�n0�����d6}��D��f���ԳZ�D��'>��w4�`}�?���IϘ��Iǟn
��_��Nc�tI����3uqK����� ���cEd�t[�v\wb�%�Rj�%�K���EF�zל}f��DaA9�x��QκA�D�F��K�v���2s�]�,�L�b�9Z\ff���畲���>[%
@;�1�^*m4�9w���M�t�����ir���'���v��+�����_�\"v�J+	��4��'���3ŝ%Y99��M�EXm�9h�~��J���H3o�
3)f���z�Du܍Sb�{�NZ��螨�(����^\#!u����͏e�+czL�����4t�r�Zzl�[KzM�.��x���ы�,��մ��2�`f���h�ˍ�Yeq�R��������Y�OY�6�F�eP�K�Zw��s����>~ ���?���"6Ӗ��CHۗ��J��_�g�Y����F���[3g��ʮh���f؝���0^U$�O�|�\�~�g'�w$�U�������<B��7��.	�:�wY2b��F)�:6���MLͫ�U��6C]�P��aϺ_�<1�D�&l/Tt\����_�a�� 
z8#g�2�o��*ϋ�N��8�}��-#ZPU��.����n}4�[�d�_K�6���K�d�4�堾�`Pޒ�jҾ���P?6T�y^�~\+Q�ju4�PkS��eK��9ê�jΤk7�3��Vq�����r귔��J_Wj~�I��yxǃ�%g�ɪ��Za�륓3[Y@����|<���ۖ	�E)�q�d�`�<_�MD�Bɚ�RX��L
�̇��#ߦ�uQ�T��΃�.��t�|6�>����NZ�3?�
��͍��q,�%;��҉n�@b'�$O@���g۪8C/�a�j�Ke-!� HƜ�����:1��~Q�N��fN��^��X�w�_�r$�AFY�lv[.Ă㍖��pU��;�bA��ZAy�9�P:]h[��"���U�G$�Ҭ'6瑚%��!�o,�aK�r(p�S����0�?:L��J��uX�6���O�D��
�.����!Q�c�q��L�a
;6ӭj�ȣ�м�7�c6<ր~�c.@�y(q۱��Z]Ô�=g�c�X<άAJ�+���2�$uD��i���L���m��e��3v����X�I��n�]�2�s������/�M�~������lZ� ��F]-l=�2�ꥃP���r�z���D�@J�'?�8Y������c��<�\��� ]�Gۋ���ǟ�+�;T'-���IC	6�G7I�Y~[��Y@��ZF�� ��=�<�9_�
@��Sپ^:�8>�i-�I�vkKx��p���N��0�*y�m���Z`����fV)is�5���u(4���i�D�ۑ�^�i1�s��c�[9����:v�[�e>�������N�OlUl�e�'��u:m5=	j��a��jV���kyu8�������SJ�UT���������,�f*�;|x��ʐ�by���M�c'{����mG0��Z":�Hת8n%���N��se�x���Y�\"��K�F��&����s�*�������n��K�8���2����M[��2<���-Gm��re�al��ۜ����ޤ4��N���2��M�oe�(lk�R�.���LL��L:�R�&�>;vDuN/hZ3�47���B�6�q�(�M��(�׹-�U���(������Y$Z(`���*]u
��m�o�V�(�ZF���^o��q�&G�Qc���_�����qi2��~��)!��S��������26�َ΋�<���r�Tv�1�����6qifӉ�<�y��7�hYu+�d͐�1OArA�\���.+����j���ű��{������e����N�-���]�2Z9dA�Dn-um������dx��mM�T��U���޼vy;�����q/^��l������ӽK_��x'-�QN�Y��asv�	�b`+�:�,��@ݮ��Z�{n���:Y'$[	w�������z,[X���Qo	���VF5�3Uh�r��sl�p3�W�M���l��6���!��8�R���U�,{�Sƒ[&m��Z���.d�]o�����%��T����Vi�7�$	,�W�8P4�Z��iq�?�ž�0������*P��+�G�1C����C�s�/�|��X��c<�q��r�o����ɶ	�~�,A�^�s�~� �P�w-�N>Y��G��)D��n�;V�b�6�奴4�׺cM��{p�kI�R����AT���ǂ%!ENޱ��1[ߖ��-e� �Q6���R�͸��|K�G�然�蝇m��j�w��J������}>��OW�"� �7z��l�������?;�T��g��sD�$���c{=S�+)�Ԫ����u7#���� �"4�=�a�T��}4��عE�J�s��H����|m�V�;>�]5S�.��`�Y���[�)[��[�l�c��ݡ�2���}�:B]^�lK'�1�l�����X�r-�,�������U�Ge\T��z����R��Y-q�I36����V���7�"�)��*e��������CV%)��IgO��`�.Oǖ4sE�^n����-V�m������ޱ���&�*9����q�2fת��ꔛ�
ld5g�����scQ,��i5zb2Ǵ2)&�i���	[F��Y�?�a��q/�t��Mk�t��$:������^�aJj�#�'KK�IKP���[R�hS���gڲȟ�����hLj5]���p��K�Ԝ�3[�^\��8bK�e3i1��&�� ���+iҲ.�*�x���ru���Ѡ�t��*���9<��l�0m�㐕_W&m�/H�m�~��e���o�A���Ɯü���{��M����u��W���Ǚ�R�F����2��G��^\���:�9�����ףa�i�0%��[d�Q���L��0��J�M����e�J{\�����*�8[D�)�y��֮�&�A/��u����,��8��A�������u�o�̓�r�\��lA�E3��9��L��9+�qfVL��o���ø9�l.m�b�X���]��Zb��r�)+o�-4�ߊ���F�:%[[l6긤־���T려���3u��1y�:\��Nu�E��mn�<����?{��]f܌q3X̃��<Ý,*�<�<(+�U�'�U����Q�\�V��4��V�9<i�g��wEw��`�$��$��h�6-��Z&��5W��UJT��p�,���2��5���L�*br�K�ql�y�F�^��Ɏ�3엶�[w˙T%n��t�ӱ����
�Ή�Q�k|9���gƂ����!�x�c�8�&��n�x?�\��U���g�2HI��-u�@��'��jʖ�:B ô�j>���Z��6Yj�^Fz̋R:[&B&���	(-���yM�*���{���.n^>���y<�>a�Κ6N��3c�����eV�v?���î`�'�_�qvG��*n������1�f�V�*�oki�DY][Y9�۬^�Δ�MJV��8��ai*�Ue&c��K2V��&YQF�� e`�7���017�������9]%��A�����[-�R��߂mY��V=Do^��?d�ֲ�HOF�ZG�����ˏK2|�LLkBe��-�j._��gX"�*��L(�b�R.4�[C�){�ղ��l��~ ��+Ѹ:�i�+cJ$m+o>o�g���c�D��p45��l����K�(|���E�zZI -��N�倫�� !(SO%���gf�*
 z��L�<��������x�|ފRo�tTw�I$��K�%�h�����.�t{ɹ璴d/��y0�T6�̂h��dl�.\�����)��E)	W�g�E���:���Ag�M�.#�}6n��+�B��I��Y�݉y���%�rs]��ss}�s�>N[_�,/q�I�2H	�ux�yY[qZ�XF��"U>�j6����\[-�+��m6��P��s��~Q���zM-M�-,X���fۙ�]zE?�A[B"��A�놼e�R�^�����v���2��t�(�SDc׹,`�_2R��*$&��P�̖X"���E"�IzO�Ad�XFS�9^�n�@���	"��j.�i1�F������iWA�8��:��18��7��3[��e1�Q~��t��n%�-�~����lӇ�ދ�|���q��4V�H[v}Ҫ\ҩW�z��l��ӗm;���g>w&6�K?��գ���T%�H9Eg����p��J�ud�f����P�)��P~5bˑb]@�����纈�&ұ�Z/��l�M�`���.�a�9����L�aDp�t�G�jA�;$:�߉=/�^{Kz�i�)�"f7ڢխvui��l�~z)-OL�mjo���x�uN�$1���\��9˜��M��3�U�Y`4xMZy�%�|M�����*k���F�N�k�vX�AT7��b%%�������9�U��{�� �򴎾�D����sRr����z�se42�������A��y���v��jtӠJ�����>�\�V�AO�$猝�����8A!9��.a&U�4�j^�nH�`��P����^ԁ�+݌�����?�c�"G�|F<��|��t��8�YQ
�&-������;�LT0��g���8�@Sr� �ضbW�[�Ţ�-4CU���%�[�mnQ�t��"�)�����z�Y�M:�xFs��ɬ��rV:��3�{�H�]�:#��;C��u�#�pڬ:���*�!�:��pQ��qڃ����-��lE�rleZ�t����������Ҝ.n�E��.���w�0��A�ƒ��󢌏��OT���(����D�J^��%n�n������Ro�0I��� �bYR�|G�Jl �y�U�d�y�b�G	5o��QWvb��T�R�����$Y�,w���n��>#�-n���_�����D�®��m���ǝ�:BifW���K�K�-9�+k+���im�f�:�)��%ni�`VQ+Em"}�W��z2&�p����o���:�������oZ�C!%�f^oo�(�9�y=�Y{)Q$�є��s̠���i�w?Z���)�}�nt�3Zfb9��d�c^j�w�=d�oNo%!(�e�jH4���e�WB/hA3Ⱡ�dq'6C=��*��"�ݏ\mn�7gUX�j-r9��߭"m�E�d�5������L���!��G�n��z�ά��+���)��u�F�׷�`Us;�&�<���K�{�{���y�j�S�[m��ݗB䨒��	�ì�s��z4'�7e��J9�u:ΞkwԱ7�weg5�kbci��s���6[�ߡ{[S�<��)N�)d`!=�uy��;�/�e��hl�$[�k��k�Y������H�Y���/�R̻�1�1�����k��s�fF��Љ>��54��k���i��R���͏"��HY�r�r�m��ױse 䕒n $��{q��z�4Z�vG{��B�Z��WlO�\[C�� ���A��S��T>j7�3Fʼ!h��0�<�i
P�:g^��!J�|�2��Y��:��b�9�"�S?�C�#��+Idcg�b����q���IkG��Ύ2۶j�
�qG	���i�K*�L�Q�lJ2Z-�^$ P���uD�r@�~B6���R�&���F�s��o�5���}����|���+^���駟~������|�_����3�s�7��"I��b�-F��j�����/O=�����w�=~�}e^V���0�z�K^��RK-�첋.�(���{ｗ�?��Z���T���Hb��P��
+�@�/~�_���޿��o=��}������1���\gg{�(�����-�d��EY��'��ԏ<�Æhu����֦��n��/��P�a��e/����Eď�� Q�T��@V��/})#��!1��n����kJ��Z�&�UJb�R1����V����^&��
|r��w�!�J���fJ�<x���)@~�h���<��cp���5]n-a�����Xf�e�Xb	�O�t{��������W���\�3`����J��vz8�xř9��ϺIꕯ�B5��7؆Ž뮻�)1m+:��A[�@�+_�Jzf��h�U�:�ns�W/��)�w���:�41;�5l��VJFc)�״nn���	J�դ:��{%�/���#����ӧ���6,%d�gt܎��	41L?6�ٝv�U����̂_Xk(�D�p����{�)�� ��"�_k��薹��Ofg*�k]m�1������C�<&��t7������e��Y����]�T��G����)=Ct��F?U��f��Fk��j2f:g����霕E��K����\AJc���9���&tҹn>�u褞���RT��� A����9Ԇ���k�%�g��
s�G�)3f�gAaH�˰a�?���,+��Ei5�P����}����-����]�,��[P5�,��3
.t�1�B���ФCVV�@~Q��H��U6���t���,ʹ�u��o�!c �7x�J��M�_�ũ�G���B��`}!�����Y�e2�(�'�3��_�k�!�x����uC�Y�-P�6�#$�aÓhNd�n��D;Q��/=MN�pʏ5��O�	�aM��04�2���-:\o��!Ԗoa)��XM�Ű%���<�*]9Q.�\�ʒ(I[u�Uw�u�w�*@G�,�����p�G\t�Ee�Ű��O�`n���_��׾�����pl�駟~ꩧ�9�}���֊X$�ն�r�}��G �~?�E`N8�s�=#ԋk�4�U��i�Zy�w�y�׽�u�Y]<�X~�e����g�}6��=�9!�5�l���{���o�w�Lg�w�y�s��V 쮭����?ӄt������,���Z�z����N��;:��l���V�J+��w�eF:��y/t��[N:�$F����b=���P�>��ַ��HK�e��t�\q��ƙ3ybsP�d
;��O3�mn&���+�9��/�<o����2�M6�d�����1o����Ѣd/����;��^�~��\"��W� ��e��Se>����rʙg�����/�l���m�5�XV�~���7�=�$ ;�Fȱ�n^�r.�j����w�k�m��۵��d �p��hb�SO�87��J��0{�����ax�/�r���/!`���LK5iy�<{@� �@X�������o�[�XNd���q%�4 ����m뭷��*0	�4j����������o=��=zq+}��b�
�qn�����K/������կ~����_ƵM�hAFh��m�ݶ�v�EY�J�O1���o��fYq�h�ٶ���k�nGB������⊼	��ɝwމ�@��-;�a��4J�k��0����W�J��A��n��&V�׿�5z>�?'��#�%b�P�5�yr��ce{Q�]�*H(����2�q����3�����W�AA�7�/�%�/=H�u���,���_��6ZQ����b�,(���%1��$}�ﾈ��(�#�^x�Ls�v&\�Q=#�eA����W���TI���Xٟ���(�v�;�w2��\���v:��*f�m��$ݮ�ڂ�H|L�	 ���툒<=�\#�!eeˤ[;;�/ �ѽo~�!�֪�/�裏��⋁L&iE�ǅ+�Nl +b���n;t;$��{9�n�:�(�Yw��A.��{�嵾�oD�0�8 ���@w���`��U�@���đ��vK ��L�k���ԑҁh��~;&	�nw�Y�g�)q�����l��V��\C�g�4�r�G^r�%r��i�����H !1���'?�y�ߜ9+����&\�46�`h!��ѹ�Pˀ&�:���?���r%���F��A����~p���3*X''������Ι�z��BZ���sx;n"3²�9���#��S�+��MX�O|��\Y%���_�t��6C|��_G ��㜡h^���������#}����UVY���?���������Q����)�N���/�t�M7eF�����N�hY�C?r�K
��� +�ЇP|�l����j�Fm�������o�G��頷k.K.�$_<��PR�&�:@���'	x��A�(�F��~�!Y��$��H+��Ʋ.���L��c�������O̟t�МY��z��y�{�G>�x��� ��	���t~衇\��5Nﰗ����/����'�q�M{G|�e]g�u�����7�gj�ŕ�=���1��)�9�6r�G���C�tx_�P�Y~��i F��I�s�.��~��߆�Q���%�#/�������c)+����qt;!���ַ�j��O����!?�я��9��0)>��|��@(�H����R�n/�{W��e��:��K���	����?Ŷu[��&����K;�#�чz@�)xn����?����Q�w��d������o���� 9�M�_���'+���0��7R��2��F�0$���7�ɔH`�/������Z����.�'P�(���|���,��P FŲ��0����_�u���� zc���}�u3�[�2x��n��`P�:3�s��l�}�A�0N�iG%+�eR�Y�9���?�&��:���sBc�Ȃ�ѹNt�;�E����;��ʷ�B�z5|��
+`8`XnF)��@ǩ$	}��^�A���a\ؤg�j�i�Ǡ?��%�M?36'|  ��Ն�t���ei�Ih��|�;�gf�!��g�8�0$�#�ˉd�Ox#���8���1�X%���<��G�A�K!i9���� �����/4��/,�r��A�cd��^f�e�*n0<��A������r���à����gg����E��|�3X%ǹ�k[ϴ�T�O��b�ۧ>�)��,��w&�`��i��F�7�|s?�kL�(VlN���{�:�-��`0&��ɜt�Iw�yg� �Р��_�0���~�ӟfXΚ�v.q�q�� 4:����?>MU�G����׿�]vY$�S�F�U?U
Rj;L�Zb�`������~���n�M�8T g�:��/�K�=���7����xǁȬ���ũx �b�=��shr뭷
�S��Ɛ���g��B5�H'A2<i=�r�����}�v��t�@g[�ؒ0ni� ��4O<��2z��.	��&������xEi��L�w��$2��S���W_=m������o~3�e��͐���F`
��f5��v�Ǜ `Q �4&�$�Q7����D�!U�)�
>e�O�p���]1-�������~���<�Ӝ-�{G��F��o��4`O\�@(,��/Γ��9w]Dj����BX��]>k[���i���[n��{�E�=���a	ؾ�z\�3҉2!<ƚ"n�-O>��6a:��2(�/~�x	dp)x-��x���<�3���ݤi��u0�~��W/�{;b%V���9ԃ&��wS3^�ݪ���C�B��T�$�� U�d���/���3ibZx�Y���Q zT�"OP�9���F�5Е��}����_���v�u��M�'���(o"@�d��W^�+_�
}��z�Uݦ�//Q�I}IgJ����И��}b?9UR?QP;�J,h%K�5�;��ZP5��u�]�a/�qƗ���/�[ h�N����.� /E=��w��G}t�lM�U�z3���v6j�T��$��>YT趤:{���oAI�X��ĉ[n&��cp;���;�2ב#h����O��� OaE�宻��B�;Jv�F�(��O�*N�螫���1�*� �������" $E���7�?�(|4�cE^,����@�7G��&6�
 ü��BR{#7�����������/�|��U:��1x����[n9�l�n��3)66�0�z5zoF����f�]v�1CJ`�rh0L�@@��4��"���D��� ������O|Q �A�t�Gt���$����1���d�T~
YC�������i�g(|{%���4��"W��a.@V���rȟ��眫���A��Y(�F~����J�1y�%U�18�j��0js;'R�c�ў�!���j�־�}�&�<��#>�-ֳ��Gf�Q�,�
X`��p-`�x���w�����|q'�#�Y����A�Ӄ��j�ދBC-Sa`��(�**�F��8~^R��EY�nQO?���q���j�:�P�n�3x�PV��;ڪ@�%�:��Y�sZ�X�s�C\%US��v��Ⱥ�0����0�nBӿל��}��?���+C.��ĭ�U\i�`§�~���[����n���{e�S��Pޟi�ҁ�w�yg^����c���\hGp��n����6�jhC�!y�Gxk8'�שD?уf �ȔϿt�Aw�}�M7�4H	�U:S�t~�l�����ѻJd� ��D�=����ʯ�ʢ0S�p�iR[!�'���`\ �k
�:Ͼ(�	�dim�8�Ou$q-0�O<��%�\2���II�|���k����d�
�yA�!?7�d�P��{�b�$��	�x�{��ԋ�����ctM  ��B�n��	k5�#�[��rIZ!��}|,��n{�a��pе��r-.�	�4�؛�^\�/������O~RG�e���ê������uRY4��<��@Tl@��3q_lH5���_��T���8�\�b��&�4c������E�zqp6���1˪��A� D�9��q��f�m�p�[t.Q�FC@����9���T�r�Ճ�+��"�/G��ǣ������o�_��ycW>[���0&��Ul�9⑗�3�O��G�����Q���1]c�$a��b�7��Mx�̚��4�6�PM)s�0
Qx�%9H����?�)p3��eUlE�jB{l���4d/��g�)X)`�G��Ī���mj��rK$����Z�]��9�3���o6�Xo��k	Ă}�a����b+�c�}�ae�0vȧ�s)�|x��t�\�:���I^�C��/��"���r������n ��ȳc����"���%q�ՑW����8���vԲB�+����z
n��cW�������g�sfLU��򉁍*�L8���6�����?�c�/ϼ��� (���)���.�w��?�a�IӐ0<��so�^��&��uV_}�~���:�gh2�<�A���h����ܲ�`�}F�%\��p�6RL.���c!n���K/��J���$fhE���o�7�P)�ٺ�R�CC�!�O�J��k-B���*�3�{��,|�� ���FIx��a�Z"��@���U:�:=��ɰM��%_T��k^��2v�$L6���9��n������D	V��LL֏z;x�y����ގ�R��*�ee�U�ֿ�ZV^yel?N&��b6�?�@��Q�Q]0t衇Ύ��ŕ*����w_a����x�� �"z�ӟ.���jl'$/]����"�)r3���9����먚R�^�s�Jem-��r��dw�խ~�����g�M3Q�DO<��4+��1�t�S�j�|��g�y��N�)qb���,P�%����L���q_��@�c�=~Dk,��������D��A�i�Yt�EѐW\q�^RyJC[��D�ܯB�������s%�]vYl9TU��i�i:�K�h�<����i�c��J+�Y�������k�yQ�}Z��T��[n���/���gu��x�'��ع=1��t�m��v�G�h�������� ������5l{W��o�fW�����A�g�q0IGq��r��}ܟYk�Y��Hq���c�3�	$s�QGuϗYl��V@:!T+��[�����w�_���+��G}�Yg}n�]�7V'���Q`�Y+4G:',���$0����K7�#K����b���'�Z�VE���;<���??���T�N��p;H����Xh��xJ�Cˡ��n%�z9���A�QPFr�u��)��կ�+�ȜL�\0r��G+v?�9��� ��կ�xoR��B�����?��Q٠�fS�V3�72Xf�e��O?����g/���2ϓ�zV�e/{��w�hI��c"oᮻ��;�ض�zk(�wu��m_|��^w��'?��C���S@��dmY�7�A�#�<R~�9�2�����[��,�*���$&�駟�[����/�}%�+�b�7;~���ṽ��ȁ���~���n;���O���1K�뮻�񨿜��Kջ4�!-6�]�A	���ĕW^	���|Qv;�|h�7k�O�/�a�t
���~�њ�<�\�/���K
��6�����F��_�z]>�����E�r��n�-�t�i�eǯ��Fi�(�d��6+�
���a�9�m��v;�:�P��(
m4��޴�mP/ ]�g��f�?�=��C��"�<�s{#8-m���	�C�Q��;l�M�*��J��u�GMN<���o�]�q5�^��HZh�Vh�g���9���K�7����Ij��� ���LǞ�½XP��SNq����������,Q~�2�7�*
�{�i*��F�1�KOj]�!/ց��
����u�Y�
�U��S�)�)�y����@Z��c�9���V��"�%W���Ճ�j1��&/k,��p�9{;��� 5.&�Q�iVcu�*ܾ�曃�; ��r�-�Va[Y���r����n������|�nѢs��k�!OەR:�� ����W:�AWQ����Zk�tV�W���X�q���6�yȮD�٦Ʌ�%���^���Yd*��t��'�8����&6��6�l���=�:��X�]l�,O�� �q��Q��G}�"�Y��c���p[��x�p5��&�J�3X�lI�	��_�r@ d��B�e��+���lS4��n�^@TR��m��h!�J�֬3|Mn���i�"�c�Ywl<j��)�����oݮ�����\�_�,
l�\v�i���^�H���xB�\sM^撊�-�a%\ox�H�q���đat�_���\$F}����]��ߏ:􊋃t��_�ɶ^`�&�Q\L���%�oI���q��ft�'�	r�4z�L���Q�F����:W����O{�U�'=����g�[��~�(	��"�6̥)��1�ysv|)��KHb���ZH�@�ee ������)��|��G�Ic��Px�Lu>�de=ރ��d�5׼��KM73��D��6>�^� OJ;���$�/��Ր#V֎�����������-o�ѵ�a�s�.�5[=�XVF򆓏;�����:s�zq�OGS�b�X�izV#Gb�dt:։a��q�1���Ћ&��LΎ;�m�v��]�t����n!�_��%�~���.I���t�sE��!.+@�A~3�7�Ƭz�e�)��0�03�>?j~gH�Q���\5=Kl����"&j��SO���[�����N����:�x��G�"�(��'|��sϝ8;�.�0�햣q<QŕOU�*�2 t:�*9�ُ*m��p���zq=���_!��C��׿��W��-���ֺ뮻�Kz/��֑���^�t��'�2��>ǩȺ���t����;�C%�2_Y�[l1�
��U�?3�Tѵ1�}�UVA�^x�%]9q<��Ȭ�ߏ[:������{|�y�M{^H�5�M�;py/���I\A����yKD�u̎��a�S�e=�j2t�n?��3�j�]��ɌP��;E&v^ŉ8y��?����q�����..p��ĮrLV�,�f�m��jg"ԑtT��
+���:��`00�I'���O�[��4��0I*>1����Li4ON�a���ۧ�6#cZ"Ǹ�t�	ҏs���n4�<01�0o�-ừ���k�@q�h�j8��|��A��t�������a�i��0����W�
O(��V��{io�N{�Ek��T����V��Kg*N~����>��c�9��=�*�Ȁ�<f䧣�e����3`�[n�ވi^ELq�)��5ȴȐ�}	ԋ̨���0�4۔��݆A�}e�5GX�~�QG��ߐc� �e��N��xK?.$~�^��V^y������4=�z1�r��L��r��1� ��l�	`�d�u�]�>�J���Y�5�rk�ѳ�~���K3/.�sA�n���*�=��c �~W�qKPG��`-ͦ�����i�M �/|�}��{�8� u�����[�٭jR0UE.c��(K���I�U��>���KٷZ�o7�iGB�`������qih�u���C0��ī��mG��^2TF��j�]v�e�hQ�iTE�A�~��M�F�ǯ_DL�'�w����.���Ye���P�G1��T����cI�&������[����2z�z�~���D��txO֑�Oh��2�r����ʠ���N;�4������,��\�h��V�-
�ꫯ��:ē�SL��B�.�L::��@4X�2�RY_�.��Mx��DM��e���->)�F4S�I!�7��NfB�����o~S�����+�^|��Qe&Kw��#d�|�u�EM��3A�6�.��y�)8#Ku����VIx�=z@��C���mG�l������+1'�]W��a*v4�,)4��Gy������c^�nbH��,��zq�w�cL��vf�nd�\����9h���j �#�'UE�������E������ �,m�����7:.�\�i����M�>���cW���?ѨY��0��{b�i�37ɲ'�²ωK�,obzf�Q:��&��R�^�kZ{�8^����im�j֬=~�]wݕ�ɐ�������|5��z���h�\?р+����rK�;���ई�.;"�1C�-T�$�]�9�����`P|�ɜ�~��8⭀Y�(�@E����]�Ҙ�2�|~����3]� �58S.д�j���V���)I	�*^���(<5������<�:n�X�iu�tsb����22�*�.���} V�oW�D�����a���V�I��d��������bQ�*i���_5��2�.�3��:����J��'��3�l
Hw�JyT�>�$;J(M��᪻��6��@�gMG���U*�0�!�B6%v��T��AΤ3�z���p�0N�Y��3!�0�I����0j��+	ך�=�^sx	%��O�m�^JIei^��������b��}.og�ʸ	I�`tZ��Y	���Q=�]����9x&WG������v�m�����~��NC��0*a+a]N�'h��r�$�"�9�q4~�M̮��a	uNR����8i��J��<#�f�2'��1�!`A���R�'�Se+e�Z{�ӈ#Q}qӀ�YI��x�H�R�XFG�^~CXr���h��k���ނ�E맒ҁp�٩"��k���u�ם�
ǋ�დ���U�LE��I�n�o�&��� �?��3��P3�:���.N�S�Z�-̄%d��]6�}�x2�"�Uz��M��^���-�d�9��@��rCӞ�g[5k�ii�"cⶻ��L�RzNU��K�#!�}4��림�K�YϖN�_�$-����>�V������2&f��T�#�n���ɲ��W���Џ;���l�Њ�n"��Ւ���j*9�ώ��0e��V3�u�R��p�k�E��,鰲<{�����f�,���QIG��[�D^���69vK�qS5uĻ������g��猵�!1~VV�$Gs�L���0�-�M�^}2�J�}d����8�M�"���a�a��S%�^\�PRE���)�HyU�~���z}2��tH�3rj�ev����R.S6��ĭ���(q�f�]GU�;dv�?L忴�Z\�*KCj��c	��:���7�K Y%�W�K�@�q�C���̱uSg�4���Xhº�@���t�"%�r����>�Ɵ�qlCϢ�D+,-j�41�E#9��G��֩|Si��\�θ�[C��8�jw�s���wх����n!?��!%ѳqb�xJ\9�Y�R5-�!�,߂n5YK�����45a�ATh�"&��B"x?U,-��9zî�k�t��QЩ��c���(N ��Mkn�����~T2�-s��c/���6C�+{��-���2Gޮ��mwe,���(������������
���x���݇Q�O���;�&\4�"��r�����"��cW��p�|�U'Z�=oj
���V30}��YcYGݦ�H�>���e��A)�ܵ�r�{N��@p���GK�!��O�������S7[^/=,��h�vuUor��B��aH��^��j�ƭ����ֱ���0��֒����_E�X?�7�m�4��N8&�[��5�ѝ���M�aT63�^��Nʀ�|�Io�L��P3��n������@�ԛ3ӷJ�uAy�F��ŏ��?���g�A���QԀ�=s�i�
t�u��nސkd�8ǆ{�-HضLjo�LFRF�wKx_9���?��CZ�ޤ�>%�\����J�X(cd=���n��j�愤b����M�<0��ծ2Z�h��A���@���U�ЀU��5��%B�9bb��a�["�q��C}ǂ�@�jh��(���P	,�~_iY;�:m&�bH�gf\u���o�wػ:���'�}ꩧ���ng�;��Su+�L���nT)�Vb^{�zF�qe�V;\/�=�Z�|�U�Ep�.:,��x��MY(^}:�VO�ל�\eG=��2a3qO�j�w��A��gK�*���h��R(�J����"³�+'�����1�x�Sq�lp�7����L>���^E:��R�a�D�*��:��O�,��t6��qwu7������]�����nK����������&�7#�(u�w�*��g>%
�u�]U꧇N�t{�wNTU�8(Y�؜���y���_�3|��̮U���&r	[ø5�+�<�=��c�?l*���9��<��ŕqF���o��>��������,��h2�n��@��c5�RR�N�]����Mv �Rr��������y;�u"<��	�������y5Z�ڜ���s�p��u�u
6��������z����` ���΋r�ҏ�@-��Y��(��]��ͬD�f;n7:ɤ�";6�����aΜ#����'�g�)����a�GyD�KJǄ&���=SG��� ]"a׋T�h�xhH�6?n����Nf��B�p�<ЏJ��� 輤-y��yL�#+��'���yK�5�����n8V�B<fk8�j\�����^M�1VD�g)�j�>��W�\��O�����w@"���/}�l��\���u������+fD��w�q��yM�>�XOӜ�K�3zFzL"�x�_�����[�Zb&���d��m��ΔK������`Yy@ul���8wk;�y��Z�+� Y"3��H��Df/v�ݳ�Y֣é�\k���V祢��Xl���'FI��A�3k�RK-e&43x Y!g�H�H��<���	"�4� 3�}�2�uK�Z��.(@9���X�gP�|�����5�:r~�̃d�O� d:��$��yV�J���Y8S�N��6���n[�a��t]່���5�z��y ����XN+��3����uDܜ�!�A4��lQ�ТJw�V�y%>��ћCD��}-hފ,d(b����T�B]}�,R��Hq^\��e�<���ꘘ��J�����,J�-n������e��Y�_�ț�TF[a��Q�#Yx��ZN��.������jL}�߯��V�:9a���_)��P�؞i��[�Tf]tь��ն�rى������x� t�Zay;�
�j�,E��9眣�%0���1ɺ�ҫ��>~Z�m��S�o̭H'{,Z9u��o��7���)���i[+,8ۋ�f�~�7 �h�è$�'�/��K,dƕ�%N݉½&AS�⋺���]w����� ���W]uU/�e�N��.QU�ֽ�����D�)_�yW��3QP
чX�]G_����������}%t=/���,��Ȗ8G�̪��a�a�0s��G�k}w�r�-��*f��@���,2*�Z�_jW|E��$��j��/���Қ@�䑭`&�h_)�����F�X��b'�kFo`Z��������oV�G�����l�)H�A�[o�U�x�v]L~��WYe�^{��;�����6�#d���Ib�#n��:��Hv�����ē~{i��*y<��7ނc��UX6븐���P�W�����a�Pwf�L�*_
ۏ��:ߒ#���~�ע�w�K���1p?���4�*��?��`D�b�q�83Q��dm�&<l�����N{�u���^��YC(蹕&:1Mܸ_fHwLlb�믿��o}+�ˤ������_׏b� 2����8ް����k�m�f��&Q���%����*�m�%��!f�?�y�BP4m��9��#q)NS��[����HN���ݰ*�ey��XV��Rg[�_s�5�nb`�]EՄ^:n�;1`	��?��|WHi��0;�c�+J�ZO![yn�t��=d�nV�X~��Uc-W��&L��/��xX����0�S����YM��;Dҋ<3p���z�+J�dGĢ�^}��{�i~iFʰ��=��v�m�)�RRT���	����uG��l:*�!�9��7M���TwN�i&���Q��]Df�h ���V���giT�ᢋ.���>#{q���K�(��0I(X��J	�a��3���W_]e���B+a��{�yr�)����[y��g�
�6���eQ,�Ʉ?�g�ݕW^i�8��jt���n*��o�P^v6ou�i0A��b���\��3�=Z�����a�&���-T�AX"��O\ez6
�Kcj��Z(2�|5R�z�d���lS��/��r4����1Ȁ��8�7�p�#La��9�H�V�k|9D�h�685����`�W4����	�h�����LUg@�f������ݖ���$U$�
�j:K|�y��J�~J���o��V��\٬b�em��u[ܹ�J��^�,)h�;����i�s�2��3�Ɛrk�B�u�ӂɄ&�l��X]�����`jM5�z������Qb�����)�]ٗ��3T�2�y�8�`|���a�W[m��)����8D��o�[��Z�Ql1h2��<�L�R��
�K��+�vGF�*����E�j�U)1Lo�n\�7f��s	�Gh��A|�푹�L2��Y��.�l�7�"���zv�J:ͥ�8U6HYyFY�!�lc��`~��l)���K�?6��;��_�c@��_\������K�6�1_$�9�њ3��c��f�m���~�/=��"�# ��ۇ��-F�\z��/���A�IU���
|��7���ĦW@�{��%��t=0L�ju\_(�+�	��>��n�喾�L���:�����>,�݃��	 ��/~��_�ؓp�Y��{�޲��S��Y Xk��ֳi�EbX?���+�'��#ן�0dv���R��7+1=)Gq�\�ZԄ�C'�'툶H��Ųc���8�a81OΕę"�;?�+��}��\p�6�l��(h�S!:����j��Q5|q~*��5��:tc ���l:_���'iU��H�e ��;O�D�I��<����VZ�?���t�=!BA�����B�y��z��@�v��/}�N�5�쨋�P�`��_�鍯��y睷��+k��ye$`b��4.�, Jȩ��	XR���LSI�N�m�� �(��`�ݥQjb�X���K����i	}�џ��g�vX+xc�4���w�q�	't��4/�	���k/�}.�ފ��X�(*��o����{HKs����!a���O?���1����RDV��'�|2�Xy�vk�J��v���>�9��{,�<�	���r�-�s�G>�t7K�cr%nyL��7�J��|Ȧ�me���A.�n�6����q\�i3�vsZ����2)k�����?�� :�9-�Pt�P��G���i��B
�ɲ�����.� ���!4k�8�CU���9W[��� J묳�Χ�a��<��9����?�x�]���d;e 
���N��5L�
#�\�l��`�)��i�@�]v�e�5״�묳a�س��ȱ9��S�}^�Xd�O�q�}�-�P��x��(Ƞ99��C��;NIǍ�8 �~��Aձ�h�'T�����0��(3��h ���ҿV|6���sR�t�aR����q�HX���O��_��2�Hҳ4��J��u�g���d{9���S��W�Bf�Xb�j�Dh_#7**a}y ���Z�Rm�����%b2^-�h%M���"��l�[l/����L���g��s9��9���+�ĩ34���U����8��]�	�~ʾ�F�4�0�X2�w�'-�G�Q���[o@�Y�ױ?l6(�e.O?�4z��K Ѣ�-��s�%�87ɩ�"�g٧50�t�M7Փ����i�[�ֹ>�j\u�U���m�rZ ^�*�ɡj�e)�G	���(��xU���1x��g�}[l1)�k�-�Ǥ7�����ύ��c�����<���m��������s�QG�`��]}�����a�7FZ;c�_}��x��H1�"�2�!A�믿� �_�yf�ш ����0J
���4xF)���	)��܎ᘗN˔(g�`��]��?V���:�S���.���+�7!ϼ��|���o��|���]�6���_ܿ� c/�K��K/���ռT<�+Պ 3����'��Z�O3�o���n��������򗿌�W��Q��)�ChH3l��գ�Z�*s��{�g�B�H�!����8?��O���h����O���7x%>?�����ED}���ֽ}��Ǟ�M�������~���:�W�.[��$l�$��_�QK�:���_ {�{ߋiG�z��LA�VK�����"0o�/=t�I|eT�$_o�	E�(د���(*ã�һ�
�<��w��h�K�Ȏ��A�G�;Mu��hQۯ(aخ����P�[~Lpk�:%!q��>�+��a5z���1��~��/~��ӛ�
x�
��!��i��0�t�����Q���:�	(�PG�O@�T��H�뮳v��=��F,�a���h����(kŶ�Y����}�sNQ0�lB�E�+Xٯ~�����1w[Gf��4^b��k��q���O���z��Ї>$I�F[Ǟ�r����B=�����c�]e�U��v[���iO�J��
�`PJ&��.p��,P�G?�ђK.�IV�l8z�����ng�J)�%� �B0!����u��W(����z@+�1�:�,��y)˔�c��o|�(=�J��p�5Ze�P;�ӤӔ�gV4��2a0z6��M�~�fm����F�2�P�����ߑ6��*���t��6-�"'+{��w�����NH�����������ؔ�E�:����e�]����z4��)�����xi��67��#��n�X�����?��@!<��Zc�5��rKûz����\�橧�b���8�mΦ#�p�.o��=et�;�07�p�n1\�8c͏?���Ë,�H�I��ߴ�_B�aIuOm/���\!����/h��}�k���cޯ.�S�d��q>��&y���N:�w��]6�UJ�1��!�Y#�
.�N�b�'��0���j����zX�`�������)Xe�J���C=��YY��֘g"ǲ�=-���g����6�d/��r�����>`L/m��l��L-z��n/)%��
l���u�]G:��<53�����
"�.��܋ڰ�I�=�zիZ��J�M½R�7�|3�e^\�8��X��?�t�FO�8ji�KE���9�8&��0s�-���(����~�_��*��M54J�ķ��'?����ٸ�D�X�Z���f�������9k�~4>T(�OE��[�3t
V���<��Տ�w�h�#����;���+�Pul��s�^x������|�3�d�8�:�%���������ַx�c�&o��u�BϾ��/�~��KiE�"����x� z9�b\��mx�8�G��ۘ&On��&�}�I��mD5�|��+-vҳ���9��&L�R�o��/"��!b~����{)yY0j��{�[����>�CqU$��sT6|ժ��r�.�sk������!ܭㅽȎ�\xt0�"��%*!�t옯<��CLy����'����2���y]�e��-Q� ����H���J :e�u���x��ԠU19� Nf��*����O?}�����G>�Js%,�큂�z)h��Т��+�%6mXY���FEKDΪ����eA�%0<������뭷�z�-�(�[q����"]�������7;W�HN��#���K���j��v![�n� �u��r�UJ�װy M��k/�P`iA-�|\�=����ٴ(ݐH1�t{ｷoo�S��`Nv�nGi��Q��M��d���K_����;�^��c2�O>�$#�v�0v��T{0�r�UWp��8��J`�l��D9W�B<����G�E�t����ޚM'��>�l���OZwӃk��dho�_~�ߠQ��^oP�-��a0� ��t�h�y�.���`6��?�!}���g�(Y�(A4�.���iLX�/kw�!�u�Q��c]"����/2��b0�� �&�
��acL��eLC;'�	p0f�"ܮ��yQ޺�m絳��l�#����?_�'�އ5��ҫ(�O<����3p�S��F�#�p,�ֿQ5`��n���{�Ys��|ΰ��~�3q�lg}s�r�7By���J��g4�K�����Q5PɁNoj�h���g�u��c��*�f�䭀A�_s�5���7A9����y+�[a� h3;���{ ����y`��@�6U�Wh��/_�����on�䀗�-���'��� M�u9ҟ'��BM����.c�n����G}�9�,x&�
R��0�{��h�B��^J�@�����W�j9�g���zx=����oա�\���\e }*�?3�,*ZD_�s�m��?���cE�+0�\a���J�u	��_�,+��2���lI(P?L2ҢT-�܎�yQ����{���UW]�;zUQ�ɇ�a#���߮�q�/�t�$s����-D�>�y�Sz�O����w܁=�<��#��R7J��NT��_��6��R�PԐ����9�4���ĪRK��8!h؏~����k�/�.u���ˡɥ�^j$�mC�^lAu�2c���^�: �]�vb9� �\r	Obe;*��F�h!x��,�C�rك5�'��3���JB��u˙���a�(�_��~��S��(a�dB�,JFN��O�8�x���-�z|^��)i�u�ā��7:�)P��6�H"Ѓ(Џ��(,Uw�f9�/�G7�i����w傹�XX/�?�3[bGRa-.���gG���7Y��_�"\Fd��BK�[�8�ÀR��?שVc9E�O�O������ԍ�ø�R_�h���~J�q��c_��-���Θ����1�\�U�4�@x=}w��A+����G��jv*��1��H+z�����^$8թ��CY|ȷ��Qf��d��g@��ۏ?�x zOXBpfRE`�"�u#G�Ї6�tS=�KR�Gˇ���cl��z�HvTL)�ad�3 ��|��p86Lef���^x!��ui�y�6��_hu��j�w��w}Tq�I�aC�<�L��Ta�u���w2�W\Q��[��7���$���@s��P{b�a�n��1}�k^�C7�&��f��se�*�F���>��t�h�L�ˆ�w�-�@=F�P%N���n5m�Ȋ1=:����v����ʈ�3����M�Ӣ��$�"�!�"l��6��v$fӅ6 	BπqY�����d������k����7�xc	���#�2L�����^�Ӣ����Y/���j�yӯ$w�gxVY���k�u ;�-�a�����f�\ׇY�DU�+d	��w��1�OJP���YI�Q�6�d���Z��e���Y��?���>��=��ά8e?�	t������E�+��Hܧ>�)(3�B���;6�-ݲX��qWI&��2ً.�˨���(@<�r�O�!Ÿ�]t6�mo{�V[mFW�U���a�?�pH��mEoJʸs#�XTV|��a�7�h#8[�L�+w�W�Hcs�LZ/
��F/���]w�[���묒�}16��W�*owD˜<��;ꨣ������-�a� ٠1��J�9p�O�=l��3���a�����������|�v#QXb:�9�����q��)!��CI0��_�z���9=���;�N8ŧ���SSp�R��%,��&ozӛH��!�us���~��`8��o��Y�Xu� �u�A1�]w����}�.�L��7Z�����T^c�::��֝��r��믿n�!��u$W0�=/b	0�z�������S�E��.�BQ�Xc>QZ!_��Th#�W���D����aQr��`t
$B��))��W3JP��(�����;d˨p]�/�ν�:���E�пTU�(_�149���1o{�ǆn��*Y�n������ ���T�{M�_R��X}�]vYi��d�ܐ}��W8�mu�K,�G,0���f�g�I.�l�.4��SN9)�hT�~:�T��F�%b!���JVs�׆	�Z��Q��⩧��p.�0r����Ϋ�$��3b�v���f��ە�/�	�C�Y~י�AJ��&���gEf�`����^�~�9ɿ�����Nm�s�d���w�s�9���t;���W�e��>� ��(�L6=�T9���SL���z���s�H��US��O��o~����<N�Qk!	�X��v�}wt�$t&���p`FQ�p{w���Q�r�m���N;�9�Qȥ�s���c�NW�~����Q�/{��{bL{�y�aSE���t����S&�s�
O�5����b1�y���]�%bs��M7݄(�*@+=�XL���D�^�ț��-��9=�@
Tls��
�k�:vrz0�c�.����믯jN",�a�Y`����5�;�XI�&!��,�����LY�l��xSAySkE�l�K��I�|wF��c�IVV��eF�MGΘ���g�KY�fW��aCF�z�x ��P���P�NBѩ�� �P��ř{x����~��q |?�tL�Pь��8�XF����ٯ���Jax`R۳����C0�0�;�E�:�&f��V���o�z�%��m��K�'Ɣ�P�AiR��g�-��l+ĒS-a/Ɗ����^b���Ȅd5�W��c�UJv����HS�3�Ȝ�Z��+A3�)wx�^]q<k��
���&f%P%%v������(l�$�bס	��bB)SU ��)\�,��^��	���p�T\��d�=��Fzt���qΰCi��	���k�jv��u������Y�^�B�	!V !�2l��	X�`�93�k�w��+;IW��,�P]�8���8λw�q8cN�܁k�<i=��3��i�!9pGZ�͇k>2.c2I�N�h�8�f8V��\��v?`�� ���2ȺD����z�\����#�뮏\�`K���'�7�)�.�6")�@���`�^X&�@��D���++�ɮ�|];�~�����.Jn�q������AN�'����_H?{���憥f�t=�5aT?�[���]�v�ސh{�R�� �_\%��v�j߮��?~��;��q�����$���I��?qC��˗/������'�>����]Є���ĝcp;⬰=Ĩ2<D��wRZ�D�'P��|����g��yW,���.@v���In�V�����u��ͤ��C���WU�wq�^��|X5�ׯ_ݮ�/�l�c�N"G[���K�3ɔ`_��Un�|V���W�0��9����֥��6�CF��[w̬C捶ޓ&j�� ����X����T�5��l��S;Hi�v�����7��|��O�p;�kc��vU�>_���v��c�	�4�\*�DX(X^�6��|Y�q���.3!���]�rh={Z[�\ԟq7�7"S�g���~} <�s'i���������j;}����Z���&���r����z�wܭ�O�֒��T�*O�\�B�{2n��S�����An~���zl���ޝs��B����1՘H5ʍe�?�|���۷o�l�u�B�E�m�[��
��3�k�Ǐ#<�]z�i�~���Ћ�����r��w�;��_v^ `9�$�ϐ����m�1��w��[j�����6��Wy��)u��V_�]k�MU��*��^4��Ծ��%�����4q^⠂�ۑ�K=�[�L����0I��BybN$�@���9�[�d��+���1f��¯�15x���?~��u�`�Ms*Y�`y�;p��z�����Y�Ł��s1;B��v�=������ϟ�W�G��8	�M>wӫq_��'���1Φ�9�i�[���u\��v(�T��L�>�eE�W8-�vĥ���1��0���OEú�����b�$E�FwG�D��� 5XjX�A�PP��ؐ�.�݆u>.C� 2n5�s�����%-�6VO�ኋ@F��l��v���T:M�Q�ɮ�^>QȠ	��Oh��q����E�c��E�7h]��O�l�]s�V2 ������t�cc/�"��b$���:��H^h ��3��V��$^�w�U� va\>$����:s�(Ԙr�REl�=U������u_b��SI�?�����X��q��b��ݮ���H��[��ܐ�[�ND�l�4�.��i�)�h%I�"���!1�r}�('�@�p��Q/]��p�\-te�Q/)0��+�0����b��	*I}wM��J?���xr��&U�nu@P�-�m��]�����IՉ�j�s�w�|R`���4]snL�$��c�#��m�S�K����B&�E@9�d�Ӥ>�vW>邎2�c��A�����62!�KTM<��M�s�˘�Z��߻�aw9g����q��I�Z��ڛK_��I���\~�2iq $�f�?5.�ɴ��z9��p��U��"�Ė�
���G�zK�:�ԐCȖ64��w�hO�-a����_�t��9�r������[�]l�����?�;�K��+�ӹ�RJ�Iz���㢩��B��˪��0J	�8CH�+Hʨ.�mԀ����Td]�$F��'5[�C��қs�0G��R[Gж0��EI�4L�K5e���ԵvD�Zq����h8�<�Kw��wq��;Jz�r�.�֛�-,X�����^�����FW��|���F7R�:@B��d�Y�G
\>9�����LNg`W2�-|�j! 0����'w�<o��e�Ǩd78zH� �TKo��g�mʂHx�誽�6�\7��|4^Ɵ�����E*�\��Nق��#i9z���m�W3����K��Ȩ��ɟj��F�����Q�:.��'D>y����h���$�X�QFefի*���*T>J�:���W�hc�q�~r���O�W���L�v�v9bcT[W���%�����5	�Pjt�	/�M�I)�D�y�+D.�O.f�\�P�a�&+��0�\z!��Elu���ٔ�i�d���a�K�--�pՆ�5��FS��{'�e�FM�슧�Cu���(���9s<+�����j���ٮH���yC�^BQ�-9�G�]Z�.�4T�d�L�,�H�p�K:Zg��R�RG1N�؂�⿈+w7�&��M� }_�(�\�}%:�0��2���Om$`��ԉkQ>��~��'~� GD��Q1G�`�_�~��������Zl��V|�:k"6��!q5�Y�m�t3��NR���+/m����z*��dRrR��&���M��%��#5���.U�Y�Ζ<��^eٚ�W���sf�,��O��	mb$P��Ç� G�OBfYǷ�\mrgH��;���$5
H��ٮ'+}Tҭ����0�������lK��J�J�TB�t�h"R��|>b�q&ךⵃ䩲�-�X�ud}�u�>T=���u|�\��I�O��)d�?	���V�m]I��0N���_֦m)�E<�y�y��p[��"�'�e��'���!���6˩�G��R@v�o�(GT��8&���+aMTn"��DSAs�s/��^�v�A�vΈx����>}��*X��*~x�[�i�*+�X�z�/��;^U����]'M�̧���#����&]���3�Q�Ť��;��Z�/�j�
,�����i�1TK?'�@���M��E9�K�+F��wE��^9R�־�rt��F0���X���vT�Q�с\��rjb-�*=������.�P�?p�ʓ�\��/޼yc�A
\��X�3]L&���Ô<�^��Q���0�u�y����X�^�I]X(:I�nEO�흭]�Vܲ���ֱ}���'x���<}�����$t�Km{���L.
�sz�DծV�Ȯ���/�cIC�6%�[��q���
`��).A��TN��{���Rl�����ϟ?��O�<�A���.��P+�I�m�]Rs���G�5ju�O������T�pv��_l-bՉ��!�@ݓm�{W�r��v�a�d��6�BHL��#�	4�S��c�3.7��M�.�I�������v���i�,j��Z9�֥�wW6ٌ]@4�}��&r�_k�v�nk����[�_�W�� <I�Or��O�J'�'naT���=z��%w�q��E}����z�H���T��yqR�ڦ������a%ۯ'����\'A66��,��]�G����VO��t�)�G;���.��.�}B\0ʝ��6�6�K������6���.%`�`�Un�?�z6����g�y���c�ZN��/�:��1]�ۤ[��ʓ?u�$���I����/�o8�*�/-q��"K�    IEND�B`�PK
     T\�j�ؖ  �  /   images/2dd0ce04-414d-4887-acda-26c206c9abda.png�PNG

   IHDR   d      �`Ϲ   	pHYs  �  ��+  HIDATx���y������i�k)k�J�d���v�m�T�V��V*J{iUQH���(�BIQYB�=f�dI�nP�c�]��{�����c������>�^g�ԁ�?�~�5V�X1o޼;�#''�~��/�3g��;w�Ȓ%KfϞ�.]�lٲY�f��+WV�Pa�ƍ�5���6lx�g�ԯ_�q��}�Q���;묳խ[7�N�:g�qƪU���٣�k��;�9sf��?���tл��	|����R�ʟ�yꩧ:��sϭY�&8�s"r��gתU+�v�ڟ|�4� +)IUѤI�R���?>���ѣG?���C���o~�a�]�v�ƍ�ҥK@�Ν5������	&t��	L�:�gϞ�>��u�]'吏z�U�V��'�hݺ5x��'�r뭷�kp�m���{�t�~��cǎ{�����?h� ܯ_?���o߾}��Fػw�����g=z���1c�~��W_}��/��^~��K/���|饗.���+��bƌݻwoڴi��W^	^|�ū��
���͚5�B�d+V���h����:t�`AV�^�
�o��ҭY��]�vV5�W���+��2eʘ/�|�r�2e
x��קM����)Q��o$��O?i�DL�>]S����5�����'(+- � ��^_��{�?�[?:Z�v��Gٚ��Ç��#F����?�܈�ȑ#�����/���W^�`�d�ٿ�_��{�n�e˖]�v%&QT�عsge˖W_DMPPPP�ֈ��Hz���q�F$(IQ�U�mŊ%�(M@�**IQz-�!�R��~��#��αc�>��C�F�b�|�?�� ����_}��w�}w�}�f�@���7onW��7�t�}�¶l���S�[�n��r���1۴is�i��*8���%��D��\�}o�����7�|��26R�~�i�^� �p�_|A52�?^x�'��Cn:��}ȏ	�r�)|p�e�FfL[[���?�a���iL�<H���k�X@��N�	P& xca���ysdN5(]��o�̵��\����0�z	Я�uH�9�)g� �T۶mmpZ N-D�W��}��������l��C��<�e ����V�2����?o=4��9eR~*��������7��۷���G$��c�E�Ɉ�"��N:(-��)��Oτ�s;<�"�>I���+��ܒ���>?<�T�7N�X����46��p_:P��/��"l&M�ء}{.�a���_yžx��.\��!r�7���/��6\�h��O?MȊ"aC��>�|�瞎��{�naC+�K����aC`
����p�	�5i҄��%�\B�����8(�!p�:}��Q�n�����K�4̆u�fIً�A�/��U��ڴn���jWV�=_�;n|�r�͈�!?~��ך2}� "�zD�2 yp(�8s�h�7�^�dIf�={��!�Nz�"�K���`�ݙt��9�ב�5Oݹs��x��8�ڄ��� '&`Uw� Ke���"�ԯ��d����Ȍ:����?	�[QVVV!�C)�e��N�{B1ee��%_%M%F��H�:Y�'��g���%K�6=�"��6�L���.S��J�*-�$��B�Ep�܁��wԪ]��Æ����4,�»hg�7yr���?>|�Ӻ?����>��_?A��e'16�?��aC�cC��!!�E��ۺ]:?ТE�.]�:�����-l�ϟ	��̹	�i�ֳ�6�1�|���C�p�y�խSG�7i2s���ˆ�l	�6C`� 6t�s�:d�{�l��5qҬɎy#�o�9LD���+W:�ͭk7oʨZ�ӛ}V,[�����V-�.]��p�yq�Ѽ�0�w��Ȩ�����1�0��U�C���c�6l�4l������ɑ�æM����K���7�f66� �n7�[���˸/7w���O<�mά��U�Ɔ~/]���G9餓X�ΘZ�����8:9T8XH�0gqj���m%v�2SeJ�.Y�$���y䑠t�Ҁ�DJ/Y���W��	��mZ���6oٔ������T��2�j��D�>T$D�HDQa����X�J��Uj֪��q�D��۷m�W����+kVf��Ԍ�|�VI�tZ�"�d���]�L�r5k�Z�v72ݶm[�j�oFnI&	(*�d���R���0�X��u>2$lh{���o�}�K!dϝ��a����wʤ�C'��b�B_M�8�������sϱ!�� I���l����oӦ��m�s_]�ƍϺ�UK~���~)�I���ƥ4�����!�o8���q��8��w�6lx�޽z�(<O|ΤNC/-��G"E;��"v6!�K��!�����uY�W,iѢ1�g0X���E���m�<�F۾�VΝ�����[��:o����*�'P�[�[_�5̈Ar�k�M�>gy��/Gmݺ}��/�N�6��%�s>�x����$Ī��w�'�Ɲ��,��b	�..%�p��׬���w׮�.X0oѢ��_=��7n���pqw���.A�y_1f@׮]�H@bL�Ƙ�ȡ^㹹KR���rԟ��2T�Zm��ͤ�ޅ��U�j�#��u��j{��\�q��ߎ��-mQ�jժ�K��;v�p�+W���K��T:Pu��W�P񈌂ҥ�Z�~���ʩT*�ؾ}��" Dd��(2w"U�V��O��}yeJ�s�{챿��[*UL�?��CJ�˗w�g( O�J2��H���D2����w�S���3�8p��yu��!ag��~�K�ݞ�>�q���0���]��v
*�ې����m�� h��X"�%تUK�9�� `ƌ�Ml(;@��?�>������}��O?��k���Խv��GNC��;�6�9x�~�i����K`ʔ)T�q�S�6m*�4?�6��ق���/m��q^s�5�HX���t͚5#]+����j��4h�9��#��鞀�z�,�}r���P�m�Ɔ�q�����:�C}��t��#�x�Z3�Y�S�N�_�� u�1�K�.���E
1�1Zl� m�2K�p#Z{��1G�P���;w�ڵ˭�޽۾������xI�|�ʕ1�T�TISŊ+��I�bŊE�Dİ�Ȍ��6n�(�~��6l� �����[��y�����DR����J���H�XD"��ᗅ�R�v�g�1c��݆IX���mY(���@ؐ�� l�}���-����%@��tQ��������S�z�z���:�w�%�'l�NC�S6�ׯ�g������.2�fC@��>c	0��L��~"�YlX�܉���OZ:R�>țМy!Q�"z����lҩ�Tjб8x�`�WcN�j¡�#{C��k��(���^��X��� I����^�%༗v�Z�:v�x��ǋ�m�;�8AKR�zui`LV����ӧO�M���{]��Zlذ! ���-bP9-��+-���j�nԨ�(%���(rr%E�ֵ�}��Ŝ��	|	𝯘����4"%��[���>�z��% [P�~}Ƣ���C����?8�#ב#G�m�5ʌ������D�ѣG����+ "N�c�x����g1��u��t�Ё�Dڷo�]w�v�ڵmۖ�E���l(��)s9m��@�zPS��w[�n��ֻwow7G���H���܀��d�T�1L��R��ODh���uȆ2SFM���`:�f�~��D��f6E U{ mO��̚5��l��#F8�@|$��I� ތ�:�qj��"���t��%Gsh��P?@Sf��5 b����\/�I<_L�=H���M"1��PC�Q�W �)2����@Q-��n�    IEND�B`�PK
     T\,b��9F 9F /   images/1d10c801-e2f1-4174-9a9c-587482dea60d.png�PNG

   IHDR   �  X   �;)�   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx���g�diz%v�	�>���o?�nzg��p�$E���.�+H� �|� }�o�W- HX-���҃K�Ù�L��L����.�қ��q��y��FDVw�\@Q���0���1�o�o����ɟᇏn��dȂy�Y� ́< ��A���'���Cd|&Q�<��Kz�\BP)��y��>y/�����=�_��s��g��];������uO�?pׄ��o�_#���E�=D���1{j���d��H9�̏����i��k�������=�JAh�e��1ǚ��o���2��<"�ΤUCR��ǡ�{8!�2�N��g���.e�-��SO�;�{kJ�[���"Tj5�#��V�n[O�5����~ah���ЯG�����Y��i��>�4Y�\�s��?{$�'�s��r�O�%��K���D3����l��z��c��t;�Q.�E�d|�^k|��%�����>L���K���d�����#��##�[{x����\���cT��v ���$c�8ˋK��c�x0Bȁ��mXA�y��֨�Zi� ���F�X�$�v��'Gؤ�˹�v8�����HÐh�|l���!�dDJ��
�U^�ϔL8��G9�D�G��Ä��M��=�h�7-{�k��f��`��*��B�+����
��^�>���'R~��`cc��#n4��%d�G��u�1*�*�^��%��ç�c>�q�����9,�%T(h��=�� ��hh��4��Q��+�kF�S
�.�'�Y�s���V3�E�W�\���<�q3�F<Ľ��e�i2K�=�ب�s�Y�)�5���ܔ�1�Y���}�F�N0Z[w��1�~�n��0)6/hqF`��-��"��](/�C/�����О9�3-W(\S*������ F����Z#�qW8��1V�|���P۰�R!�Q�i)��=���v\� ����D�� �Bj�d3S&n�Z�i D����`���� �5�,I�¼���St�<&C�!.w�&!#2��7J�_��Z���b�hy/~G�J����z�?L����󅴙��e
�
�D�j}=�M����a�j��TJd�
ʜo�y:~|�\j׏�,�p��V�����jD-����;w���6��d���J�J�� ��ϧ�U0ܬ�;9i/H��1�N�=/�D����{f�V�����a���\�kkx�����2|LM�r�c$��R�JD5cΨ��{Q���^@�/xN�L����g�?_�z�R�y�;)�b�tQ�Ђ�ň�I�U�GYh���pƉ����/����M4��)G|=�=�偿�`	Lr�1GԐ)U��O�t�0������6�N�@��D�7��]c�A�ǒhd?_0��0�_��\��X*8K�tnng旰X��Ώ�I�!%�Q����nvvqw���?p�B�%�~Ñ��ը��0L��d��cە)#L�/�[�����ؑ[�S�Ä��u%�$���&̗�e�5����$U��d���CZE2�or��[[xq��UW��b�o?�p�u
���4̌Y�R<����A9���e�{?���<����b��n.ʅhgF(�K��r���G}7���!ο|�N�Г�Ro;\��
�f#D��5�Q8�F�]TɄ~cjJ 
���'?g�J��DH�M�͙J_f�	��Z�V�F����M
@)�
��r� Y��d��J\����=���gϐ>����7�d�L�!{)�Q�PB�9�՘�xJ/Id�׍+6p�vՃ���:�*!(!B��~N�g3��&Z����Ǣ 2���*�m��{�d��-��wξ���gqe�NGsh��dUʲk�����`����=��t�E��y�.�:���O��8&m�jL��w�x��A�Mm�4w�}����l�(mJ�,��$�\��F��EA��v����e�����F�������H,N�9�<�ڕJń���~~��ydw�н���6J�C-P�)�j<��"�cO�$� �[��/���p���C�nO��rOԹ��d5I�����*�������p��-��.bqm͈��%D���"��\	UQa���?D��`�F@�9x	��|
A:�$���(����׃⧷]�}s�Ҹ�(�fK�k��F�!�Z�n�G�Id�A�Q�H�7B��F����Q�S�Ec��@��}��4��,3*��*�p8|F[� B�fsǼ�!aQmw��!mFB���MH��1_h�U>+2C�Y�ؑ]��(�А����;�_�o\~o�_�Zmª�H+���y��k�3X�rW�?����O�nb���c�%C�H����4<�V#��֞i����9�P@���r/�
��yQs�s��ҦC
���e��_F���G��m�d�8��l3eN��OIk�y������|OL"��Y9���]��Ӎ���`��Stw(�ro"���Hh?Y��3CS@J�y��B,�4�s�Hs�>
��Dm�.�(
�5]��ؼt;�=.�S�Gf�P���7:�g��ѓ�(^�o��7���g�W�(՚ja�n�ώ9�j�s�4O��Ep��!��ћlB1�و���x���Rc��8_��ZI`M�;��4A%a$�xZh9���8ђye��U�1�PI�!1t���Oc��j�,�^Y��H8a��̙VFGȰ�$5J�:�e=�f�`��MF��
x3��'Ex)_��&O��[��㍕+�����ﭽ�e4�\C�f�Rh��J�ba���x����y�ǜ_�� �qƟ	�sV��)YK��u93
��Y��	c$K�vN
�!�m�ŕ,���p�G�܄1��bL�%����˧>c�1B)�/���w6�ϗ(e﮴p��e�^\��&��Op��������
)]<�K��l�М!zo�!�Erm$ ���z�l�<7�=2�m��r�$�gIȈDk^Q��~/��yj=�+癟w�9������fK�-��[�=��|#�����S�,פ,��
���:t�<��g�/?��ıTx��wJcqc���I��O��r�lt������Ri@�
�zl�2˝�/wNj-n�;Bo�O��țx�wp��F�Z�To:.��ݼ���;�{[�Dm�h��Hmpn��}�$�M&���0��8�E����|�".�-��t	߽�:�\{�2�2q�;b:�
��c�^e>E�R�v{ڄC7&/��$�z��*m�v��E+f�������6vSl�v8��Y9���E�o�xs�M�A����&8"گE�$�7�>,���,viRm\*b�4��I��6��r�17�@s�N"lS�&�2
?8�����|f"�P��F&+�P�1���"��b /#�f.Ԑ�S�u�Ή&�MB!�g9+s��	8�w:u������iYq�4��ZůE��d�C�/�Z���dz���+2��L��(Bd��g�c�0�	�Y�W��3�g���9�y�5a�:ۛ�1�K���cOy��9�eƔ�'���ֹ��b�T#4̭������Koq�������!J�54./����޳;h�	G�MH *nx�a���M�c�̻�2��ƞ>��7�B����9�*�\y	Kd��@&L?�~&$�E2�"i��7V���R[��i78����rQ�,��h��(�ܔ�d�&��9��RA��3�>{��i,./ckc���H|$^2uD��h#i��@2oI��?4r�α �M�󤭐�e^<�v�\ڕ���r���e�����mRxv'{�hv�^����y��Υ�SD�:�&��y�!����!��p$�ȘN3��lU��c2�p8B�ڠ��c@1]�o'YS0N�c��4�?<8�x\�=�)�2M"�I���Cp���~B�}�����z��9s E&���5s�3��g�p�W3'C!o�y�TR7v�sI#��̽r��n1C/p�������n���:s����rB�4hY�:0�"O���K�W0_�M�E���]�z=�L�7-�:�"��cB��A��o���ar�	(�n���WN]���Y�(Ac�� ��a
�%/'�8⼄F��U��Xh�Q=L�I�B{j�5����k���p��3gz�QC�SA��##�K%<{���~ ��4�y��Lc��4r�!�X�V	��N�����XN'Ž�^/��[8���`k�׈*���s�4c����<�a�6E�Bc-��F�<�����R<zO�)��Icr
�>�Op�,[�ks�]�E��}�s$��*��i�ks.S��P�Иsxef���C�]�����R��hO�c�Ia)���>+z��GT9!��0��j����8��
�i�2�=8�����Ǵ�5ʓO��1���C��⒣��y}��Ơ�~C)鼐��%��9���4�xU�0F�. �3���-Œ����\)�����<����>�e��Hb襁?B�(�j����.6�`�X�%D4�S7Lm������E�˨�M��6qm����e�w<s�$��8-#'��� ��z�q+G��)�6$�Z;�%B���}���!%��n􈟯7�X]YEF�{��뽛2��Rd�s��k�WM�� I�� �_�z��:횜Br�{S�T�	W.�,�q_\Χkt�q�7!4����	e���1/tg4�ɀ���ٯ(�A��TX�35yd%lF#���ۘ�1HZ*��$;X��<�(b��p�8i{��tKa͠�s�+WK��%�x4!29�tD��sM�]���0$��)̥��,�3�&�	�L��y��j�*4��U�}�)8�=RaF;{�WNS�V���X����=�dc���3��}�"�e֑���19��%*�'�+�����ƦfS��q�X��B
�P/�r�E� J����Aްi� �B��PP��	�N-�`m�*A�a��Zp�s�ӿ�R���S`�^�%2�5Q�y�zh6"1T(���GŐg�B5Q�:�3hȗ��r�������%~�M�,�n@F����*�YH��98@����QXR��	��DT@M��2����G�pkt@{�3��$\A2H�y��%��[h.��ݡ�帕��O�$8�FnΘ}ǥ=����Ӵ9�h(����s��eu�-�	�r���t�ת��*�@j�_�`h��|&�4<�g%�Y7r�P�����y�6wyDT�[e�	���X�x
g.���Οǳ�mn`���PGI@��r�݌j���;4@o�1�oP(���(C<��)�,���W_���K�-��������&~|g�h��Z�}����?�V���#�S�I:��q�}�p����P��mgx��8\�0'��C�;J��`��fs���G6CՅ�k�./3&qU�X��]��'�!�/�f�W�8)�X���HطT����	n�K
�Q8��}�#�1A=)�m���ְ���GP��y��'��6P�vΥ�bm����t/�@DI<W9����s�d����85�^"A���RVP���&]�.�;GH($#e�dNsX��mV`�]SxPg�M�ba'��+>�}����YKz����53�.	����e��$j	@�Tب3HH�	�G�+5b�9�f�P)g�Wנ�Lc�?b��ϑ�KȚ��p��~o]{�Cl>y�a�A2���p1'�>z;��PK���D{�+���|Xi������9�[��d�Vi�W.���a�g�O����l�i��^�cj����$n����|�ի}Jdy}\ɻ�sԹ�R��\XJ�m���\��C(Z/�m���-s�!w"��R��̊�0x�G
Ԩ=�
�+U�6\nzX��pޔ�&���[���|��X1��	��A�ԩ��xc�#+���<ơ�g)�l��W"smlP�tP���S�e��l�FsΝCx<�����ow��r-�ҞqK(c��'8��.��زQ����N�×���p��ADXj�V�{B�)r��%�
�Ϊ	��&�?7/&Lع<�<p�,q-Ħ5�c$q�ÉÁF�$t���%U(�����5w*Od����bg�ʆ��c�C5
E��aiLAC�__P���Lfii���R�'v~u"�����=���Op��5����d�[��x�B+������歴��\0�bIJ#Y�~�"M__Y����A�W?�'_�ƛ/��������
�'�wb^[)��K�ڐ�"� �Y�'X 4��x�1ڏ�a��,���~X|'s��0��B�h�v�����m!�,�<�1sW7~��K�/�+p���(U��6:�c�U�(M��Wx��8�LPx@�ݤ�M�,w�"�/
��=Is?������&˫�+/�Y�2m��#��,���S�doh�/]�DB���y��Z���h��$<j�a~��������8ߒ�=0&-����M"yE�=�!��V/�a�`���Y��d/�����-�6�v7Ao}L�E�{�� �r�|0�>&<s_0�5dR��������Į3P8B���@���x� �G5V�!���$��
����I4.I'�$��rUsg�H��q��S�����7~�\�mM����w�Γ�E˃"�.�ח�(qM�d�չ�&��+X�s�<y��u
ͣc<~�⅋(ϣE����0��5_��_��R��t�sM�q磟ᛥ�(-\��nxf��3 �QC�;�� ��w�8��T�����4pCt	�#�y�L���l���:�����`���vɀ+�S�Zp�s�W>��H�΍�߉F7��Ψ�J+�@�2Mbc�1�XRB0PP��=��R�����i�[;��g[�y��
�mh c��]�z�\�wo�ư�5�AbDJ&��븾t����Vk��M��#�&8�~���XE͜$L�f�LkL2��L��d�.��8	�*�.sL���L�&^�	s��8����g��GM6s�`Z^$�Z9\,:�x�����j.rl��

�X0g>�V�^�B}��j9g��:���~������\{�M�V3<Iɀ��W�$��uﾳ�ڀ�O\g�4���M4KD��jx����3X�m��-TdH2sf�$q!p8&.�^���xT�i��D8ܻ��Gx��w�\;k�rH�&m2�m�m������j��R�O�b}s�!I_^�d���l�bg᝛^�]v��A��^�C��T�Ê���f9��0kH&<F�e���(��p�F��!m�q�GI��Q8q8�X9��T�L�*���v���:��xV���WFܨF��d<i�{w��sl��bpy<������W��{�!���>�n�2><�8����o�E㥖�u||l�q��mg3�%N��\�$tۘz���}��\yִ
��l�&s��y��-�4�ʄJ�	Ki�Ei���Q䅄y>+�1ә%Oĳ���~�����R�\����w�B����)&�n��������JH�����J�'�*0_�b��dާ�[xq��3��P�X!��g��"�s��kO����#�������$�&�����3�e�ط�t���;/�3�?����q��Y,,.b<LХ��QX�RŦ�#s���e��#��8v���4��v�u�OB�-���S�Y������r}W�g���
�:����@%q�����z�GXo����1����������1���1Ⴢ�26KQ��D�\��Z�7p�6�ݍnjUe/�;ͅ���@[��}]^?�,�Ҟ�nf�	C��wct�)�C~NMiX��r��T�=d3���QX���n�GM9$��F���N��y���/��9���u�dnvTz�H�t����Dk1���������+��cB)�̼���jz�ӣ\�iFWp�#$%Fd�R�b�RpT悮#��c._#	��#i=E(Q�y�j��;zj>=�B�}>���ԩU��x�d1�f��L��{��*��G�.��/�wn-��Ӌ��P�<�ss�)�ۘo������]����	�4wP?/|yP0��-��L(T�U�]�j�Fc����!YI_z�#J��A�-$R��%�a�J%�E��EڔM�'�i���Ͻ�{���2�G�>t/���Ks����b����v�S�5'n^�+����ϩ�>r���B%SW�DU��}��J����huŕ�e,��P��x;Vq�r,C��+46���ۏ����q-���Μf����g��>\�<�)�J�6���$�4oR�+0�t<a>���c�����P��+���|f��E	�C�/s��_�*'�ډ��IƓV�]�Y0��Ya�a~�N��V��b�.e�FԠWG�T=2�iCBu��L��C��a8����3y�]���gm���w5C�v���?��M\=����Ҿu�ؑ^B=�C9����l�>n�ʿ���f?���2ݏ�9�*�QU3Dx;�E����Yʵ\<P�Eڪ��=���ťdR�<B�������"�LB),ö^��q�̍�j� ���I�;� ���'����Lb���DE�������Z�����N��
��$FK�X��e�#��z�p��>{���;]B��e�Z���*����b�?��VW���E^_�./Hs܀�7���ʅ�.ܼ�������(�S8ks���}̏�G�]�Qӿ"�O<�dΚ*I*3{ٔE�Mjl�W?&�j�x�Ѭ-���
<�}ew��]ew��xtR�a��bLS�K/�S�q|�ܣ}�6�S��rk�D�T�������)}Y b�Wt��ב����F�͓����M���ƕ+�q�8])XXd����*�%S������}��*�|�[���eܸt�7񃛏p��!������\��C��iT�mBɏ�(I��W	�*���q�����4�娊fc�3����hAjR{ء
�l��~\�]3�p;��ˍ���|�A�_�ԍ'�=��Ɓٗ����>x����"}#ƍ�+hEu�v5��̭R1K{�A���������c|�l���ͪv�g:e2�j�zj��J��"�h�T�����ζ��~�0�GM/w��ET�nO�=�X�4����/O(ת��)�7 !pcZ�&�d�ŉ|ߔ��H����N���MpMPR�7�&v�D�ӗ�/�Zg�HC���Rjp.Tm��Ƒ%K��WCL��5�f�	�s�C�1��c�{Ak�ȍQ�Ζ[9�0�(Da���]G��#oh)>���<gb��w}V
�+�zM���]X0��$&���2�=<��&�X�k�Mz��uiz�&sJ��3���;�x��p�{G��-
�Q�����*��h��x��;qi�V=�G<�y�����I`�q���2� �j�� \2Y�*��`� �H�*4P�� VǴ�km���&�6j�bY՘�d�e.gRź�I�Mn�$���ZF�R�g�=�&<�?����^<wW�`.�Z ���j��������_�����g�`}��c��!�-VR�,��P!�m=~�^�'&̎b'Ie)!8�F������b%ƙ�ӆ
޺�~��$�%N{|�R"§����}pܧ4&�Uu�'Ns��:I:�*�Nxw)���86;Hq�^�gp?5���rC���i|�q$~�gS�%RXՈ�N�l��`\4�X�;�9xȰ��
�o���$itl/;��,��R�9�r���S����^WQ�5p�idA��k��c��9��A(��foR�H[�)p�5F�i� t4�z���)���O�\3��pG+��K܏:�smm�8{2��?��7?��n�2���W��Ƿ�y���ܦۺ��R�]Ն�S�Wf�<�sPmTƽ.o����R��Va�zg
���D*��~�X���������u	S*��#@�x7u�+�C�>��z�0�����Q��;�4���R�h��'[����sx��e�]X&�$������S��|�l��z���]̉g��)VV�Ī�������"�`R�"�p�ju��P�,�
�>�}ǲ�+�&�1&�"t	�6�=�Y͜��
d��,����%'�OAx"��Z6��#A� h%7�ʤ��	'PR8��S��ג$��i��:�B�<�i��#sZX�����K��s�\'ƪ%I�G��*+�N|XA����CN*�����d�3�5Q�g�Y�l��K��Gǹ�?X���Ș,􂥈?��#ُyf�T�:�a��
�.�j͐��緶�Y���R#_�-�*��ꈊ�y��c�qh�R�%Z���(y�_�$���w��E
&�}��I�-͠rs��)'�d$�tH�&7L�!u���7�ܱ�0+ɷbG߶M�����@"�8�6��訏�oc���R%%ul��n= �m�� �w�iqb�W����̍�U:��� j֠I���PU�u\U��������D�R�7H264�g�R<<v�ȑ3o�C-p:�˼+��pLk"�d8NPi!��hhڢ+M�>6�)�OH�H�}xF�6���V<�얌�Cb
pQ�O%�PLQ�Q$f�xM��AθHҞ(#*��&�/��:���y�%_���z�	5��,�@���3������~P���ż<�J�T�.�O��"5��ƪ1%힞���|�5���K��&�Q�Z4�Z�vґs)���К�'-0�30bpv���kH����<�E�l�TE�>�l�e�ߒ=���q��c�jy��IPTie~��`�=y��+Ң�����]OW^I�po��4�:�9H�ZAe�Y�@	QH �@(�*X;�f|txh�����N�(�����U`�lз���\��j�f��8��L�aWn0�,�"��4����T�'�qZ	�_�c��=�_jԀgϝ3U��lAiV١]Z����*tUُ�xƾ�]�(���u>DUC�d8C��95���B/(r�5��	�|���W8�J`N��0J,,��#�&>kh��FPn.��9I�_�(l���\���Ԗ9���В���1VDh~��9,�ֽq�KU
<ک�c�)L��Ώ��*(�y"�P�sō��0U:������L�\�o���V��Qqk~�VNcQD~_��#Rģ�gV��~��<�7�+ɗv�GV�V6�`�2-�q�+R�/�Kibȸ�쮞Tb^���� 7�<k�rɈ�rD|���V���.�]���."j��:ڑ�
Pm*�3���>-�H��H��k��T��ò����,��}��4�}f�|�b_��ܠ���Ѿ
zxm'���n�y��hq\A[!���I:X�{<a4W�	���$\���R����1wf6��c��
$s�0J��h�ܠv2���RC�h�'q2���b���d�4ƶ��PH�*��U�+�s�v�%�hn,�����N.ZOy�e�9gK���x�Å��1���r/I�Kq�����(�8;v,ڨbLz�I+��x�d����_A��f��E����/Ą��b͝P;!�rDo�������V�;; ��㗉���ys�ښ��6��ݍG�ԤaK��(gP!<K�xX"B(�$uC��F��qm�������4a���2��,�b$p��+�^�>񹸰�&���/0��qfa	g�V1�[Dr!A@��PA��v�̹�S��9KR�\�E Nh�|� Ә0�9f�^L�Z�̟��Ndt�$\%���D��k�w������.�������K���'9[m�4,<�J{h�괎 c��V\ $S�KI�>>Y��۫aA����1����#�&e��59�*�jz'�����T�����i�'P�����l��W=dGpY�E�"������\&{�YjYFh�to7�>��'���{`sk�u���\�f��o�[�;�[6y����X|���UO=�������5K�@=8�9Bu��ū&9ZT`�5�X��c�����.j��U���S�+p�(e�C���q������C�5�}%_�T4��cBٖ"L�=�t
�D�̵�P�m��B}����%�x�Ϟ�N&\�f����E&�M*���錱?�H�<�e�1I���ޔ���8�+���d��5f��������^3���ą�-R�#m�o�����ⳏ?��;7���A�,~��t�^����Z�N����R	|��u��sH�����&�mV��E�m�R��>����Q�0p��2x����s�.�2N2[�$��&H?�y���U�j���4Lci�ܐ�a8깪w/\�#;	ٸ�CFe΃��O��}��8�q	��gN/(����*��=���wr0��ҭ8�T:!_9:\<�86�Nf�qKT����J���t�wqD#�ӧ�4m��|z	�d���m߈�=��5��]�jj�<u��V��ϵ��s՘��N�}R7'.����(���;3�7��q��F	������}5�/+C��V9���i�ް�㍎��\h̹���%�3��E�9<H�c�,�#,��a�T哪��7|��g9����}��S�\>��'(����]�[�&Y[;�.ao{G��Ԙ�U	s��J������x��Wq�Ƌ�@#�����q�z��Ǆ�;�y"������狆%�[�p`6ʔ\>�U�#+�+xJ!���3��� �o�Y͚�7���bҜ ��P�.A~B�}����{���.r/K���Í���Q�qi�=��R���.x��S�B����Q��a\5?�¥j�UW�(pm�Y��,g^
�+�[���q���\��w/^�KK�V���#K	��;ħ���@��ճ���=ܾ��l�f��B����^���V��ScdRE��A4Wo��Gut4�q�f�e�(c�~�v�ף�H��� J�,�P6��T>j�ؕ��W��VW!e��Ƭ����SVB_6��w9�9��j��(������w-~�07g�::��������ѨX
�`" �Dcm�P40�s�iF�F��]C�O	^����^��(�������l����Q2kk��ֽD��VW�W^}���_�M����s�0--��{������?����^b0+MC�|��Q9���i�B�¶ʂ*�Vg��ht�۷6q@!.s��7�Ā���Ɇ٫��uR�&c���%�k/2�|y�O�G�T��-ӻ���C��!�I��� �������K����>"��5m����\�%�D�xz(N��.J���e�~<�>�&{>))��Wv���	?T�^YZ���;��j�[�������5�9��E�:���+o��!�h�����<��%��K��9&}
c�%W��sX$^_;�s��R(�x�$D�"`�x{�n���CɃI����'�4Z�iM�q�T�,���Xo�q�u	S�L�0c>,c�2�7/�@fib}�4ۻ��Z�QW�{F�3T���Q�2�t��o�?�3/���'� i4L���O���rsɴ\ط�[�Po�|R�$j����/���Fd�to&s�P��c���4�U�"P���lit�CETal��R�$�
����eͷ�vȊ��8{�,���|֌��މ���$��&V��X����#�)p�����L���8$�I3�a�=���,���S�,�Zm���'��얀��;�^��][�c�*ar������x�睁�xj�y�!�_�s���"[̻U ~b�U��º�mJd�'�7���Kx{~�������e��'AQ�[��R�`��*�EU=����޺D�����qO�~a� ��[mV[�x�W����]��˯�,��(���Ӈ�X�&����G��_l`�P6���X]9����e\�z;�ml��PR���W�i�*�?��3��z��d@h�[o�o\����o����k�Т�W��������qp�M&|�g�y���.T��ҋ��o�������x��G8'"+�w�{��GV�z�����ϑ4c�3	�{�"9<��ZF�c���Fa3�d���`�ƙ �'T̐�3�oz��'�Q�����]�L��!�"��rR͓=��y^8�d��������]��`�AA8�i��^����U�S�>�	�Rf�8j)!M-g�bsV	����43,�J(Zۉ�ه�Ȳs���5����x�1��<��T�Zuy3`rX��Ïc�@˦�N��e���}P��7n\��.���'��_�饫��K����Jǆ�x��γ/0�%l�POu���*^8��G�v�b�Dd����W�O�7�{�k�C���8ǂ�b�2�3+�|��V7�6��R���2�]|��5j�>:�ǘ_X�2�qx�n��~���?�����P�_�~��?�g����<	s�j��N_�K���y�����DE}��J��[�f��L��ځ+��ʄy޼|�Z�-?8w����Xŀ9�
	��5ʌ��T�cL��K��=d��϶S��GQ�]�C��e��A$9C20J�)��%�8o�4g�`� ��?�>�y����\�5��jѽ,��c��W)�%L8og��)��I�Wl��-ګ=��ƹ���>*y�t*۠�%���/�����V�]�g��_�X�L��?�_�p�kg��"�����QJc�v�2޾|	���@�Ze��x�[�M�q�m�z�C�4��y���6?����%�0�&E�����ts�ٱ����dT��W_�˪�sJ$�F�{�0��v��mtW�|��Q{�KC�D�����4#����WɀC�����N.���3�����-�4�Ej��N���e.4P��S�̛Q_",:sz��<� �b��,�|i?&4[��@�kК��?v8��pQpma�r艕)���B2�*�МI#�;�;�-(Έ�Ţ����`�������0�okn!
�w���0������
F]�Se=�y��̹u����m��n�~r���嬊�q����(y"ɦ�L�^3�ܰ�9y��1��j3
,�)�W{W>�s!��Slmo�~a�R�K�O�?@�@V_��!|8x]�lx+(/���݉Qv�ڼ��{n	ݡ��S���{A�I3��>�p��+���M�3C��q��0I�+A/�^���6����z7����1m~,$#��@�T_�t���3J�\�qg� ���Ң6k��S�*%��!�Y�9�sB�*
�+�������б��ZS�̂�u��� ���1Uޤ��Q��-�_��2���qu�4�,.�SK#���};P�UHb�̩��#L��s1������ǖ�&����z2ئ��rZH���6r)�����Y(Eh_���%ե�*�U���%!;{ĕn	��sM��VG�����b��%W��x�]\0�D��ȵ�;:8 �m�7�6 >�ĝ����Kȶ�Zh�E}X�S��cm4�v��ݻ�1$��j͉G[��kݢn0��p�S�|����gz<�Nʼ}��l����+ƙ3)]O��k8S�ǘ�du�"��չ�\<� V�*�*3�B�k(/�Cx�O��F3r����.ʱ27���e�3lw�,�z�������.�[����+I-���F��:GV����9���U d�A��r�rx��kx�ŗ�Ž�h������ړ��i��<����5�(��pwr�{����$�r��N
1�0�F���c̗(�3������ ��W��9��9�EA����2��':y�>W\��D�����&�df2���
p��f�-EN��� /��Dw^�x2.R[Haoc�6��d>K��\�ͤ��d~Ӈ�f�9���M�:�G-.LDV�.���>��Q�Ba0���!ƨ��F��I|1���%��ޓ�)��.U�d��i�ua���*ƞݳ�0B�3�׉{70�	]��|^in�1�Z$�m�*���UJ�����}G�;|��S��)w2��RG�N{pq��֑u]��Ti|W(m�u�	Wv�����Ekw���4��W1�a��	V\��(אƕ����kvB�*�-�a�Ŕ�����]��m�2Uo�$����R��f��!��Y��H0[$�r(�y��nј�qhAy;|�{��=8��H$g�l&w3(ڴO=��Õ��+����Sk=�b�·?��4�Ҟ�M�9�ʦ\�nY�]�X��	E��9�D�\�^����AL�~ř�$`�-���7��o�Z��'x������i,��E����Q>_�sl��"�3g6�g���}�Ft�ݾ��F���ՈX��)�9X���5������>�z��s��Ἕy�\�m��`�:S�>�a���,-�"���	�
�Z$P��rhɧ�A�(D�W��x]��l�W���A���m�h{,���5�@�Ϭ�^D�?�:�p�A�6B�â�H��-%��|/��y����]�+oz�̂��pws��?vz]����� �y+'Q�b�.A�F2�K�ꈩ�;�^G������^�*R�n�IM3����O��=�H�
a���ɤ�w�Gv"Pf-�"rn�s	H��U�O��"�h�h~��|�l��Z\U}ZҐ�њ�e��-�kZM*�m�W�u�����Q#s^1A��`�V��
��\χ�o���w��r�������*��ؠ`�/a��+X��M�`��;��1v^R
!t;ǁ{�>>B��e�6�� ��F5�"��=�)�Z��pJᳺ��&�k
�X9��	1Ø��=jT�����f� �����#s��(#��ʓ���e
��f�C�_f�iuEOԁ�i���>jܬ��.��&.^
-�9��V%�Z�	7�h׀�����,%���t1����#_��'��b~&�v�q�#d�[��AUu,;�[pR��Ha��g�iI5����VJ�If䮵�`���6�)�j�g���=�M{
�6�7�cx<��𸣚>��0�D�PZ^�K��(hZ�'�ʢ�X�x�������攸���0�Y*yQ�o	��
ͅm$�:�!�n�_��o{�j�Z����_U|�w���k�}
ŅFd����.��j4�5����n~jy����Yr��j������ϰ��C��7m�Ϟ�B"\2�Ɛ�����꛿D�eO���t�*?TH9��|�q��:�[�^_��+��^��}`�W�`�﹵I|{��&BEj�?r����R�b�iϚ봣�PL����=�ЊW3�Д�j���hL�~�<�y��;��D�u�7m�eG�
w����Scƴ���dK^SF�̽�y���R�������;_�^7������O~�3�_l=>/���ک������P�.K������{�[��Dg�bn~	W.]�勗��9><�Fx��w�m<���]>�f��2=2�~�{��YP�������G���k-�uz�+/}��7��]?��c���1ݯX��:�d��Wږɡ|���y��f��� 17V�M�UP�p"L�`B��4<����+2b�#/��~}�M�_�n�׷Pi}����@ͨ��A̼�}8lwQ�}���~OI���a�Y��M����&T�d�D���y�Ƌ�k5��ݿ���!�1$��{��t
��\[}������$����>�Fv�M�پ2�7Y/�g��ޜ�KJ@Pz����X��5�B �����a��rLܘ~'V�;>'@4��>e>�:7�^��Qz���ã�.� v�6�Y/��[Z�hBǃ��4���oН-v�Z:�&��p�ź�f�O!����[������67���k7Ч���9��[���)7�����J]8DKvd��_��_��_���������V�Z�/]ō+�L�|��M���]��G _�Q����._�t�,����m��ܢ=*�~�>>�u��3��+�!!n�p	�+�����(��#\]���{wn�/~�Qy���gx����[%_W����h��uX�U�Y<�Zm�b���LW��dv�4�w=Tݠ42=�B�.U���[�����	�X�U��jn%ϫ�j2r�b
�@ukC��i��>I[�@�@����%�|��^u	�5
����1�ǟ~���o�7��������G���?�;�Rm��o����5��G?���w1����B�~�9��A�?f�a��p���)��܅3v�Jf��];�`�+�s��N�mk�������"�B���c>��.�{� �����s$�]��n��OǸ�Ư!\��o5����85����_P�m�������ٳM����j�h<��M��NȖ[��/������4i[�!�9�f��ܛ����ϕՊ��Dk�Ϭc��'��ο��Ў�dg�	/EJ?xp����I8�����@a��.����|�쑅
�n�lY�Gs-�G�{F�|\�:�ϟ=�������rf���)��9�ӽ]
-���<������.aY;���8�rW��î�9��G8��}��|I�a�3�	����'.�1BiR1�r���>�Q�j�Bk�pp�}��M�H�!PvG$VS'B+;�a0t��hm�F/1�'��=$<A��#���[��u�h	��!!�
�V5������C<������go���������̩�Z/AkylU�1�}�ꣀ�m
W׋��չ�y��5�%*P�?��?�A��_��J[�KW6	�t��?�`������<��#��ʾ��s��C��S��mB��.�8�D3좽w?��u\|�X=wٜ2W�����t�m�����G[8�K ��WP���QL�4��Q;D�%��A�4%� 
}�o;�D]���l�Щ�Yy����?� y�l�:Q_~���L����ˢ����i轖�P��vn���U�:�(iG����[�}����8��A@f�P�������.r�������e������[{v�W@{B�j��HȦ'��X�g"6A�ٲWo�k|��TZ�%U��Nk��V3">�0Q輛j`�c��c�Q�b�*�q�'��<�08y"mQKW0���t�
\ՠJ^�11�a�������
CBP��)	Y�V�v�o�/��/�d}�[y�EM�T����s<_:T��hY�N���|�<���h��s�ս�v������8��u��t��,�M�Q-O��v�`���zrғ(���Ǝ�"^�gXJ��x���C)���p�\�b����&�m}J�����6kesJTt5�u�7�&jcsDܜ���Ĝ2v���U�*�`xy��b���N@��"w@�R�j��?ه�52tfy�r��=V/�lZ£�_uD�B����ǅ�0p�b�� �����r�
����|��3��v�u��
���5Bse	gW�PQ�?BIi�����R��н���7���`�N�qN��u�+���ܱ/\-\�ɉ���PiqK���C^=u����ą!���Qsݞu����Υ�#EجE_dU���Q/Z##���*v���7�.���M���wr�0R6���1��eOi�.���br�����G���]�X�kx��غ3k�ʗ���r��5ε���6rU�"�3p{��R���H_��Y}�))��q��z���񰍰��ڱ�yqJ����_�.�t���Dyue#���&��}į_�k+��S	*�Y`)>svրʂ$1�9��a	O�(�~8J͓�<F%Q%������������]�Nّ5rv��픩��@yU~R*��j�ZW�2J��Y�
H�H��h6��#ߒo7`
.t��}�x�v�%M�NSu��������&�!�\������:꫙����$�6a��!�w�!gY�K�^�vaA�D�j�;����;�s8�!�`��o#��ʂ۾M�F���bU���O����Z�-�<�\O!�ǖ�U5����OK�֏+n?�&o�,8]8f�p�Z	.G����:6�^��^~�lL�i�:lDy�e�i��) e��aj�&��s�����d�Yx���4_q��e�`*��U����Y5Q��\`����la�{��?�9N�x	+Wϣ2��1���Y49�gzb�WE(��+�f:J)6�S�U�%ˈ?�x��Q��}�,^;w���զ%�����{x��������6v�KX�d��Eh����2�@q�z�T�2R�����Bb�-�2��j}@�J����sx��:�Z	������ƨ��\Nn����ܜe��s�T���!��z�Q/��,�=j���܊K�̯a���|��ý}ڤC;w�sH+��Wn`��!�.m��x�j����g/3G���VH�%��,��̱T��uwnB�s�rR1y$�S�@c�i�)�|�VT
[}�a����^�S�V���%z��FU����5UfWyO��q[�U7��tڂܲ�
%���WmT�*�x@Β�}��B�)�W��/��o�����?��n����Q6m0t���8�*m�%���x��o`a~���sǡ�6��Tc��Hl��U��J�(*�c�D��ӵ���W�;O�楴�̎1���Z����#��sX^X���Ǧ)���o��.M���{FW���]��Qv=������}��%���b�q����O���$��\�i�������m�Etǈ�ś(A�sLi6�q�c�x���E4Μ����Nb�,%U�V.k%pɦ�8�h��E\i���z���ua�m��n��߻�9��ڜ�+��cie����c|�y����XK��~��x��wyA�amB�L��q��,.�`k{�<�{��|�	�F=t�P�C����祄��g8����T��Y7wg�5i�d��m�SZ���.\��30�9��m��l���w���+�p��E|�j��"nQ������ɧ
ܵ�R-S�+�'��9�߉,6Fv(�
�`��:M�ը͑��_�3W�2B�Nƈ��ѧN��3��~�մ���¢%A���}?����g79ǡ���4�/�t����C=¿�?��s>W�\��Ԃ1�����]
�.�Qj�e����;t����n
E�·>�Pz�5)N]_i�4L-ĺ�YD�$?t�����k�v����#��Gv����k�K��p��E�h]G�I�t�ƥK�n��~�L~lv�C>�lN-��M�.sÎ)$K\lFp�O�ѡ�W�?�&/�-���Nse%��d7QE�%D�͑XX\�%� ]w��2�}�%�]:Yj��ev-I�եe��w�ŷ_U�4�NU�H���-9,�!�A�?������*���o�G��;"ۭ_`�p}�V�]CTn`�>��*���<u�E��v�d�����ؖ�ۺsqʴ-�?@�g�֌�d�7����3���6B�1�n�5�6�����s����]��o�&N�vh�th;����/���\�L' �p���RUܽs�6��_�[7�+�a껞9(("��a3y��1���Ck��x��p$"2	�q�[PYG��Nsna	K���QL� ��)iݝ�����Ԏp���Jm�tpl�TA�\�^���_�.���;�o�O?���'�q���e�?�ƶ�L�M�Uke��܏�F�Ƽ��,A�2�
ǔoD+-'�[�ݑdec��eJe������\���l�$L9�e
��������[�?��?���ɟ����8:@/Jq�r
��/��4�e%J��;Q^w�ZH�`ܗB
_�|)����Itր���"D]@�2�K�.�	�ơ��dwɨ��CJ���A�D�b	��ʑ�	�j'靻Vr��$?�o7/(�:E�[���r�}B�.|���zdj7H	~���J��TC����W�TWq0&��/�µ����}j~	��9����y4�橹�x��1~���|>���!CU� j%W��DW���V>�Z�����I�܃�C��|�R����?�w���`�B��H�]I}2���5�v��!A�٤�Gm�ȗ�1�Twgg��.`�~��]� �Z���R��^�u�Ը_j�����=W�%2�bG��߾�?��U�Q�q�ư��i?"jU�-�@�wn8�ǹ�Х9��v���3Wf�׼�h9^hH�6fX]�q��S%FҸv�Y�NRR͢�Y�Y���d�ϒ��pP�~�8��ګ������[oY���=T�bL��s�>��~�)�:����Ż��=�Kj������-��U�$*�=xv�p3��S�օOMvG��0H'n��Ǳ�p;3�֖�bڑ2�}�?k\$'�b>u~zL-�<@ey���I���댋��Y���!�S�Y:�6U�t'j�j��q���
%Έ�+�B�d�_`.~�VTr��ֳCY�R�R��t`g\�Z\�|v}k��Z1���	��H�R�S:5	1�Ң���ÓVn��`M��%�J��
S��vm�ԝ�@�#B�1?���]�p��`�$���3.zG�j�++g����U|덷ͱs��ϱH-�ҋ/,����]$8�4|9����������]#����aooo;�/�u�fC��p���N
����� 1��w�؆U�3�]D��#iڢ���?��b��+rF�lm�Y�@Mw_1��7Rpg`��	��v����,�&�4�w>�u����:��شh���iF�yT�;V���bwЋ� C޸q���~���V�����)�|���?{o�1ߺs-*����������?8<��Q����6���+��8_�r���=�C�L�n�g¯�>�2��S�*=Fffޓ�Zx'�g1��*���hp�*�I	����F�N	C��u���&��9�G:�k�>��.�8��������j�=7zw�Ĥ"p�B���UɌu2��(�y�J�"��%Kn.�j���9ݪMSv��"���32��rK$��E������fp�G}c���1�.���O����K��,"�:�v�j�ʋe\�vň�ڛ�'&�Tz�`��	�~�����{��AO�*AXP}B���F
I����se��(�lF%V����i��7E*l�������P�w��<��vs_w��:\n�53r�p;�R��d^��
��F2Ш�����SogcdEkFw���CU���4��x�A�36�E5�k�k��|o���ʕ�����m|G]�Ca�o�/�l�	��ְB�{����T��Gs=v���~���������=�w��?�ޫI����礷����� A�9C�&tG>�(BG����̓.CCr&��# @�h�]U]�g��y��Z�w2�����HTWwU�1���V�7��ۄ*��`Zv5�kB���ұl�N�s����c_�x��g�$ê'���o���(�m�IM����&��L]��T�1�02��a0Vkȗ��3�D���ϊ�gG�<���\�5i��K�n]�$�	/nzs�y��]�������lhYIFG���� ��|4�j��L�'^
�[��-�?�Ca�̠q����JGC�Q��!��^��Դ������di���D�.xeennV��&ͮ��YB��p�̥C5Xax
L�t��(��HC 5�N��D�e�I�O�n˶����|�V��v�ڷ�Cn� ?i�l�1]�Gx��Z�E��g]L�:�M�	�B�(v��E��R��cz�3���� h'�"��{���f�+"���9}z��捯ݠ�3��fa�I�����f-6@5T<�2����o~S޿���ʫ����z\��~��·�X�L�q���Ger #G�U1��q̊p�??���.�~ye
���O�k�pc���_�1��a�ow|�t���<'U�]*��)c8���/��#U��֮[��i%T�90��l#���!d��_m�B�+a:��{���A�zYC@�T�]�6��=�r�F5h���4��#(bsbp����НW���KHCT���pLT)���sg/p�==�5�ͩ���!����������m��!H+c�4��3r���Fr��
烜�r��Q��XNĬ}�G@�\��P�x>"E�D� �z����AJ<׶4� jvv���p��~���R`"���1sG��;O)ph"�m��_�2�������rB�V6=f�q͝qY҈�'�Wr��uy�"�)5���V�WaH�!�X,B���-����`:�������[�~�;�ѰWn��P�Ǒ����h"&#�錦&����~ K��A)@nM������	e��$n�Z�PSf4���d%�x�����Q�CU��J]J-�!)�i���{��X�2D�k�X
Y�p�B����H 	�P�ܚ}a8F�+�ݟ(�(����������:WQҮK,�4�����R`��i�u�o)"\�x�T���6�?��Xr���W�7(�ӿ�o�xQ�^���b�<�$D
KT��!��I$I���ԩ�9�X{"o���̙3TB(P+�ss��O�<a��x:�[Ճ�D�+v 7J�x�@9QZ�s�F$(8���a>s��]@������5���ǖ�=L[x��A��J�LA����tAu2B�l6��E=r�,k1�k$B\ݍ��8�D��V{��%��O"ן�N�6�6X\����s"�TMr������>���O����3��{����~_Ӕ���{�P��8%�΁4#-��LI[�����|�o'Z�����jN�Q7{�Ҹ�h�m��^�6�������+r}zD��:��0[	%��+{��Z��k���cՏ:�(����3�4������PƳF� �N�����2�����qqr�2�tlq�������}�O`�*$!�%�a�L茦�!�?�� �h%�����������ߧ՘<���������}�hx�N�fHW��Ɠ"��j���j��2�\���LO�ˡ�!˪����L�zTH1S�f�Q��e�0.CL�,������1�A�
w��00,Ë�r�HcȬ�x���{�|��}�'��.��%Q]�g�'�Ņ���޳w����`�H��:�5��kٚ�U�HVF�9�@���w/^�$K��9����cl�44Bk4k�}CA�t��ʹ* ��m���Z�����s�ܳ�˭�n��ξ��J4��K��X�)尡F���|�W�UCUt�R�7HN�e.��ԥ���)I�S�`ҡ�Lg�������pV�ʿ�\���K��t�lo&�7R��ɔ���&d�g�h���#_/�&貌;�����X�^X��FX�I�g��:�����*��i.@;��+�br'��Z�g6��M�`,ۡ��q7R�F��OO�AR(e  a�ԛ�O$}ǜ#xQ��G��J�B�PP���=���0y4�n���S�r��ʃ���!Vhq'+�^W�;v�t�*�0��Y��2�
��A���rJ䗖���]��H��ܽ��s��N�5��s덡`�jä*}�F��6IXo��ʨ�z��g��k��p�^�ln���d�i^����Fk����tfv���k���s���q� [糡�k������;)���ݛle4�ӄ�^�@ �OZ�y�/|�;��j�ت��NG&�俻xY�=2$�㇚H��R����G�'kJ�ܖ�fG�qzAb��{R��ђԠd̓f%˂\Q]1�-�b
���Uא�|���*.�`�����]�k��,�&�@|i�)^S��)S���۴�'Ö0�5�[K�G����̌\8�!�2>�f,���>i�M�\��-U>T�Q�6�+��\�{{{���7�y#�B���u�?;�N7Wg��uZFpC&/���㽘#�6��׿�y@�a ���t7�;?eÝ �l�L��`�];�zg=q�G@ka�AߒM�v2�ye���F�<7�|��4�i�r��9�p44�D� �����=��/%���/dMC}(��W������|TJij��b��z���Z-C���/���#��5YPK%��cD@iXԜ�ioSp��>q��m���b#��$Th���OH��C9�9�rrBf.|]�������|C
[RZ{ �Қ��C9;��?~NnQ>Q�X��g�k��,}�H;g��~)V+���i�Ü�*%iMW�	��bL7��
{;��HW�* �v'X��J�!�*
:�!�Y�H+Y���`G6����˨z7�3t����3;6��ā�B!N-����a�D�H"���!����1;m���P��;:ʱ�ʄb
�XbS����F(	hY�24�;��������@�LA�{��'�G���%V����^9uPeX�99�_�U� aWҐ
3A�8�?���!�?d��7�{�cƏzh~�j�(ulu��d�X�������!�7M��l��j^���o�y�В�'�GOfogG��g�L=y�H��V4��	R.,~yp��#?������ <͆޷�ن�>)�P>p�^�zU�~wNv���ӞD��si^3��M]x���f��b��q.����ۑ��9�>1%�Ɔ4����������/5��rP@������29:+��)l��fM.L�%aZ6�~$�� �BZ�2�W�e�Mv�UXË��w�Rh����Cy����kE��2�p����ի��j��9�ݶ"�dc���
)��Ò�)bTۏ�$=8,ss�rn!.	UĎ�M	������9��YQ�Ц�5ņ#���UJ�����%���j^��t���ޮ���{����>�$?�я�������Y�g ��\8��9�����2�F�5Y�pLU�~�z��|�<~ђc��[qᥤ�C�� ����u�7d�T�8K7dơ�f�
H�"��4��\������	�֬7��0���`�魏tmʈ�䚆���{��ڊ(����$��ϤR溅���zK���~^����]�K >�<af��X���;����65�Xc?g���@��򳂅��p
�L����j)�~H�_���)�y(�����%�̢
c�R��Q*L��'%4�ɦ�a�$�rN.��5��:���VKH�� ������;:������ں�m9*�$��?�PZ*��3���K/�E��؈<Y~ ���ܹ�	��E�Cp�F&$;8ƶC$��NL�k.,.��G�H~��ԅ�y|�'N�fFu�`ӆC]�[����௭>��<;:A����栭�,��H���ӡA�1�-�P0x^���<V��z�����Q��06�[�3�����7퇆i�x��Zd��F��E����1�bR=��HP$��,�F����[vm�E3��F�����F�*_�%��h��m���ls�����*�z2��!_VL����֍�y�\�
���x C�S�Ih$�>��ϝ;�ŏ��Ƨg�^�'ja�����z��-QGe�`Pϫ�-�u�5^'u�׊1�����f�no�jR�Z��锆rUu��3g$��������I톆�>zKIM.��9�|�"�����QK���K4�_��r3G\���ba]UY�
��G܂K̉Z�^{G6���Ră���ݽc�,�կ��4�)8�XeW��yZ+l�C�#�pYn��<�(��'�[������`\�Jl��]^�,�4�Ba�435-���9;��ٓ�w5���619Ae���W.�{T�2*��.^�n�7�|�Jg����4h%�:�O��f�J��F������|�;���;���KU�MX �B�9v�l&f�N��JH_|��H����N���:���z�m۠�?���Ƞ
��D��`����,xB[Ĭ�f1�c�k��%�{559�
)�����9���Z;n�x�o~��"����M��8я�f�{r��*��s�Y�v��{�Rji��P�Gxo���S� @��T�pK�&�S�Xt:��鸺��!It`Uܶ
^Ԕ���>c@!I�j��	�*c'Ғ���&�59n���r�Ċ*���� �2bj7����Z&T�~[4ˑ6�*�S ᠟��U=Unw_v�6� ��R�&��0���dx��b_7
X(����=�#<�+馡k�u�C��5Wm��M�hx�`ܥѴ �ݡ ����)u�4T+��ʕ"�k�*=)hҟP��N�w@�y���"��6�ՠ�>5/K�OI*���=ztxP�vAi�g�&$����dU�p\KX�p�	a,֫1����g!L,`(�[����H¥6�d��î5� �����a��?Ǵ5:��}��?�m@�3c���AX���τla���ʹ:�+�~ǈ0��෻-!���u�LMM1F�� \FU2��h�<��V���P�"�����ۆ�!�mR����=<������:��#	?,�df��_�C B�q�Q��
�/�l���#�_�j"ӈ
Ks-��rc)�����P֤�eLu�_�@k�vZwπ�AH��{���� G�����,7V#�����)��Ro7��B�%�i���谤��4�i
���[�æ��~�k�^�`�Cas�!ha?&�v�;$�y�`�������C\} �|�=8\v����,�Xp����|�S�����r���(4w3T���1Mh�9'J�y�<2XxN��_��ɤA���9�/�	y`�d�]B��>L��C����5��}�
]���T���/ XM��Y��ȶ�n���/ E��ΖX%F�z'�FBf����)E��,���^i?4��Y�a�-a�R�}�T�{_a>��^ Vp�c�&@c2w Q����͛�H��#q�{�&;��&}a��rX���Zi�t9u룑���X6*Mj�؜�+���$��D$�Np���>ۉ~�N<�@�T8Y���D�
�7�%mx#2�p�&�����K�%Ώ�#	a�����k�RF�6�j"��SúbT�TP�U����^1U���QvM��#���ך�P$�0���@�W���	���nߑ��\8�(�#��ɝ�2<:,��^#3���c5�PfJ��P84��\�*7n��ʩ��e%��@#��N}6���׺�
���yq�Fzp`����
'��&�#p���q���c��p�g��J��Y�����G��:O�-���@�c�����s��S��OMM2���@�C�*;�k�9/�̘����8&J�Ѷ3}�K��W@��� �J��-�Ԕ����00�����fF1/>�E��kQ��x�4c�#2�I��o���b	�P	��|��������>�Wڱ}8�:z�;zs���Jss]J��2q�3;"�ܟ�b=�C���ܰ`�޹-��`�( �r���Ǣ
�^��ܸ���Zu[J��=�|쭏>�ۏVe ��?����~�#iꃉi�+d���Qa���or�ǥs�����k�z>X7��� �}��e= ��@���.-;�L�1�|�� ��p%vd�F}S=�/�!�Myw�H�RE&�󌫐@XJ��9vԫ2Ի��^�����hX B��KK����U �x !kw��̦��U�WV��c�p"�E�%{ `�`�H�mP)ͷ��o���CI���&���(�C�n�. >�:��8�o����L˝ۆ\B���2?0k�hHл�|�2�J�L�2C�2s�u��ч��{�����b��l��,�ʎ�g4�QU�u�}њy��>��@�����N@�|,����Ɔ��[o�
�ci�Lr67"�g�jm�>�!�mC5u��|*�B����j_BN�У�=��҇�b���>|W&/�"^h�3mH*C�vuL�4�(�K��+-��Wdes[Jz��S���c&�y(�"�q�I_�rY���eqt�-�`�z�^�D(.k�۲83+W�.�X<#Gޡ'�\	v��9wjI*zCl>�������ol������bqI6����&��#�6@j~4L<j"�����cڴjaC�j�H@sĈdа6��VH�+4(%=WLb�R����m��{��g���T�6,��k���p��8���� ��Pq������z�
`�
G�a���&9/M#>AŃ"C��F��ȱ`�1�6���!�����v�E��L}����	S�ᑐ��U�ƁSUO:::��
!��g*\ߟ�'F6(???�o��UxU����B���fs�A�G�7==��F�:~�t����跽��;�����da~��<ƻ�<�5�ā���3�J	Ec�Po^S�H�M5����� ��>����Iɥc%�NJMϡ�+HK#��1�۫\,�M�gC���#�D^���J]`U���І���$������I�X����''�	k;�uG��[�Z���;����/��iͳ����RB����Lƕ}8@r�:�ͭ�u��PgtbB�Ge0��ax'�����nK[�ɉ1U�	�&T0���*tG�Ks������-)�@��a�T�?�0T��� |���!��$�(t��x��x"��cJ�����|Ů�#�D)�t㣲��ܹ{�Ȉ��yV+^��r5��x P�W�B�:�$Q.� BP��.��ݕO4;T%6�ј@,�si�X�d������h j�:�t!C���)���"�̈́c-��y-<G��-��<�ׯ�8�Y̓a�`h@nl��yWj8�AB�kw��J'��gw������j�k��Ny��7(�L����3�:���t�n����q��=KxOΐwG0u�!-��y��X�0�ƹ#���Ӓ�}�<k�ya�cK��V��]������F=Ժ�ݺ<>>����Rz^���x�$��Uv(���HhT�z"B��z�${OV�r�%��#��/��u�4��5��y<`'�;iH٩���0�=l�QI�������.�q!�ȇ�bG�^d&��sj5�*�Y��gf��}M������pw��{��9��P�B%�j�ba
:z�Vn5���O��q|U��Y��O���~����'�y�Zln��V����<��u�X	*�������H��.x�x�I9�tN���U��	���r_�x��G��?�������[�OFl,��6��ƩpX�ɦ�Fxn �M�9P��ƖU� �
M���}~�ҁ�����^��;�,�ڂ�ٸ�+j��rT�Q4�Ҝ4�L<��bK <�90����Xk�g��Ԯ���r���9P�����<��ӧdbb\���O�����e/���Xe��_�h�,�gA��4��V�X\�>�7�|C�/�p^�~�����ѐ*�#�e,c�пZ�^c�B��8����0�Ϸ[��u[fTN�ԋ��EZYRA ��e���V%;��{�ֱ���
c+6���+9?*�������+k�Q�6�.���ج����Ф^�Kh8�
?�J���Q����?���T(�4�f�\DC�L2i؆!�p�X���;�U��/c�N��B�4����;��+�%I{�^�s|�Uf�E.L�h��癛ر6?,TE�"M�_����Z)���w42�<vf��u�T LJ{��?�yr1T wTaQH��>=6��f���K����������z"��+CP��/��ׄ��ǴF J�0�B�>�<�B�����O	�d����������b@�ـ�'��FQ�"�biF�KU�b�e�[!_79mo��aT���Ν;@��a���S�NɥKy��݁~ �5o��6	����!|��X>���x*�V��V�_�|9��eDn(��ؚl�����I�(�ɨ�3P��R/QM��#�P��LI��z�X-��n5�uT�TgX�FdO��A]�В�BC�kȇ
_[cC&AF�<��yS"apM����L�~�z��V.*�VE��JjxB?~�q4hx}��s����c��/��I���i)k(���#���[,o��@�=�#;�O�*!r��ޅ��O��;�AIK<P�+����4Qϕ�&Bd���ZF�~�
g�-��j�Z	���>����m����^���g4�wI���5w�����$( �C ҙ�u�M\E��k�j�?�}��@v ��&�	��h������B[�ô�|�@�kh;���'���R�<c��{�u.'�A$�^��J��:��r#N�Koj�S/ ?�]�CG4�E��A��&����2<8r�Lz��WEAH	�o��z�#��*�wU}!��k���tF�67������hp������,Q���φ�Zn@��Y^y(�z��+�j�k�tQMa�TV�~C6���T��M\*[�N��[�w���+`{~�<��|��g�\��e��ۖ5������dwW��x����SɈfG���@%z����{�<�/H��#�p���Ih�.�s}"�E�b(�UC[��߽�;Ɇ|Y��`>��%[Sk���a�cU��n~ ����l��k�қ
�*��h^�4��/KA�j\C�	����n����ctԺ:ظ������5I�}�V��j��Bq���f��!.����p��S�sG����RRŪ�P$�ۜY<M� ���x�����r��!Z��2==�&��KO���*yGQ�(�E�(�)TW�^a(X~Tf_���]�Ĺ�V?j�Vt�Y��M'���sP.H��@Ժ蓎����K��׃�C`0Ձ�,*�Y�q*@#��'�WC�<�Jk��x7Ϝ>����nj({@��A%���t�!
L�-�w�i�4F���������5���S��;*;��HT�$uF�tBڕ�ʴGg㑥ϴ���vǶ���x�ky�p������7(������\Q��A��H��VX�$ʍ��]_�*Q��c�a2�Q0��~O ���FǑ��<�<�d��9��YP�Q%��巯�)��p��Ė��o�.Rzs0R�|�H��BX�5d�����32|I��̀��NH�"�UΈa�	��I7���i\!��gi���%2sgb-{�-HK��kJ|lH�^U�Ge�E�ۻ�D���+���Qk:<2"������ے+�������Lqo�>"�peyE65� �v db�4wlY���&�cP�Th9����eDA!�Jj��h4l��\��՜li�a-;��G�yA�D�cX`�����<\��q�-H��ᝯV
�\��{D�RPK�Zv��(�=X�~ݠ*��ԤTj�kJt�Q�E����w��a
b�M�����܂���0�h��,�̼d���<�BC�s����0��gkmO6�%�qehn^�5�Z/8�j�����˵.��}��,�Pw�����^�@V*(������a]=�zݗm� I�����؀T�@o��4`�c�x� ��;��C�aN/@�;��s1�o(m�ml���U�u��zܕu�������ڃ��Ґ��으�ꫲ��+��.Qh���Ұa��#�-z2}������{�=V<԰�I�Y=\�Y���ؒ��kXWOO"m��@�p�7/ ��&�#��'�k��Y�"�i$p���s�<+W5��{S��-����={�k,fh0T?YY%��P���&�U= 
.%V���;��+%�f�+�玖 sUD���,��zz����yT.V15�@E�ƞZ�^#_ț�~7/lI���)/����V��	B��a��������۶�~V1��I�yLSYxN��(��o������c~�ZBۓ����-�Ͽdo4h��):�r<�a;-�;�@x�8��j�*���ܠ���>��N����1�����IYi��]�c��,�n񫥑Jզ���K�՛q\;&^òIu@�zW�������P.�p4z�*��o�Y��!0̎9ąz��dH��&����$jY�`P\AxK�j^��������7�!X� �#.wi�reY�ݓ'���^�={*�B�l5���&ˠ� �XV�~]v��	TF�}�N�CU%��G���H��7οC���(�FH=��y��*�J�U��_�yK>Y]!j�' ��f�%
�)>���#�5��0��Z�a&Fe �j�Uc��Q�<��/��j2a��i[.K��sn���*3�Z���ES}�j�����h�M�����-`ڷ��`�B�f�FE!��>O�5BɡTXN�F~*U�6 �'@���I��z>`����!=&�KÏ�&h�'�����?��u��R5�Af���+%�cN̓m�ͪ�����'Qt5�����̠FU	�gb���gelrRr����UiB� "p+�g����������0<�uy�����G���-��n�Y8`5��+Pv���-Z�Xߵ�R���$�an����BY���-���RP
�Eð�������D��J��w�Mhp����0���Z���z��1\�U�v4` (�k򘢿UA>ԇ�5Ѥ�����]�̦��Y��d����4Ĕ�[���?�+>���S�4�p���>�u���[}ãN�*Ij��a����ڶB���F�
g���05��=��wl��K�ٶ�M|E^�B�nǄ�Au�;P��b�޼kB���������ė�o���1+�^��Td�ڦ� ��ёQz~T,o߹M�z0�����#
+�H���Lk���g.l*�j��Fet8�a��KB�i"*ە��ܨ�I!W�FN��>̬6���&*�8�j��`^�/�e$���y�zg��1��یx�!�61�o�Y{�D�A�&�骳��Fł������%p`��!�z|�GȊ5c.��N�ڠ�͠��L�3G��ɜ��>p��� "AG��=;�f�s���Zu��rU`é,�o�:	����WA�mn���h�t>�_;���"�V���[��g$T�
� �l�@��f�Q$���q:����1e�Q����I�z�:�=��0����%_e��?�280�P��n/�<�u�0�	r�V���G������阴�"����ah� J�i{;�
�mB�����:OC�fR�yڪ�gh�c̗_~�Z4�.�8�~P2�OV,����#_�l��,��*=��I}nqU�r�U�p��Ґrӗ�����efR1u
n8f�B���k}z}��~�j�ݛf_��Y
i[`gO�ZǼ�����m#�t�M��}f��8ʫ�Y��3���X�I)�԰e����p#F�s��
kHǄ�3���
^c�*�rQ�dC�Q�,L�P��unYuT�P嘇*�R��כ�|snj�d���А���Nd�Y���K0��;l&�[v�N]�=�VI�ǿ� U�
�������B5C4$����hر!US��HxJl��%�g||�a(<��ĔY;2�?����64��c��򑶥�g�����U>� ��W>l���Tlq�0.c�cl��K��O���x�����s��K`:��e���yG���v(x:[6ʨ�M@CW�Q`����C��u]����~S���T�q��Q�%e~zT�y̓5�x��#RFq�5��Ų:�fwm�����RX>�f���j�QCC1k�����c3ѯ�L�	����P�ӛ�0z�t�j͐KE�,��K"D�8$iZM�yj��n��C���}���h���G�9����0g��Y!nD2�Aa#�?؞[�*����P��CiY��������%b�NR�;&4vŬ��'��(��"�ƽ!�����B4������#��Ɂ�H|@#	6x[�(�� Eܮ�����c]�p�z��}6��dѿ�`�e�[)�b��IȡB6׆ ��{jC�޶��R��@(�?���Ì�	�!@�t<3:��쁧%�rJ�fp���A�P\��a�:6�����-�� ���!�
-���BLs��cAL��ݝ-b?S��&����3è9�z/,�� �пCH��4�>����}�M5�}T�h��2e����3���W���8�M N���Ҹ�h�����&�P8�?�&T��VϐG,ޛ�5
"x3 I0��A�@�X��&y02�s��C�"j�k(G�4 %p�A���U� ��/n�lHB��"g$in�����GI���w�pLZo�
���9�Q����q~Tȫ����a�V��nh+X�)����r�ް�&����B.��I�^�L�IbPad�&�>��F����N���5�4.F��c#��M�a��a�G=�*_�5$��Yphy��{:��b����ȯiA������Sgv���xn{�@���w�nVZ�
,����E���vr��7d��%8 �ě&\��#BHn3�a��H��%�2�1�كۀ��#�1�	�Z,Z;�y��O3d#bS��]���ޫ(f>Cr�nh.Zc�grdRBMOr����	A���GZ�����	w4bB���6�0��2 {C$��|��5]�& ���F_\���vE^���hC�4xB@!����澼�pC4�$����*A�m^�sB�Z��B>S60Y"���ox�CP�C�
�� ����(�aeۄ��*
�,�1���"�WÙG��|@x8U!&�1f����x�Mn�_y��� i��F����n�c��s�i��L[@��{�BF�B��� �SC-큾wJ�ґ��S��!U��\:p#�;��zA��k4���y������-�yS�����{����ɂp.x�� ���.�����Lu�c+�DT��1���)�I3���w�N�O5�f-�5@=��<�\�~6(���=�4��S�L��6F�RH�䮵����$��h�X�jSܲ��-S�O�Cgh< Y���^�7n�b��[o��/�(+;�`ݟ��Y��T�i�V"���/<#y��L녦��gh�����Q�p�\А��k�ƃUY��$�"��e��NZ ��E�L�HLC��Aޤ�"v�±%l��M2m�)j�1������HXe���5rIL���T5�.`M���b'�`���ݝ���E����e���1({(�БT�{��i�"?x��s;O�9Aá��j+	��>=�"��h,��R�kWk;30&cj�+��)V-���w69C�	��J���8v��M�䵃�rC���2�1�vq���aw������y�QJ�⃡��`�k�o��M�Z٤���|��`���j��3���"-�}�D{�D�\S ��wO*_�z;�l@��w 
:�9!`��y�^E������h�}��v6��AլW�r4�T�� Y�"�>�À�<iZC��̐��Y��g/�L2+��]q*rztJ.�����Ȃ��ΎOrZKX�_p�HG-r����S����7�/K�Ɏī-�����>��5er,.W�c�^�P�%�?ڗ����dW=�A����t�=��֪����4~�n�l�ҁT
��!�@��x����h�[���$��ǉa�h�����Z2.�PAHc��6��;�N�h��T����hh�4� ?�����e|���4D�%���`2{�,ߢ�������<�2��p��q�[�2�kl~^�7��Ĺ�#*�� ��Tv�M����3n���0x�Y��2w���1l�n�T�W�4�:�r�:sĶٚ��\����;;��J�!0��n<����3������kw�dB�W�����P�S�N�z�D<���Kz�-+�Ƭ��?JI����jj��D��R��҉8234%y��ZZ����4����dDe�Te
3� ��o~�Y\8�m�� ׏�V������L�O���A�����"�0{�d�þ�~�\j:�o�=+?ZZ��C�ohr*jUԥ�ZzQ��_Pa��|{M���:5�J�ͪ�k�|sY��(C�=�+��Sf�-1�d��D_�EUE	���������aM�q'v�xj q�چ�<�Fe<��%��<�BM^�x�}"���X�l��\?;�wwv�w��&�}xS���V9'���m}�~�就��@SS��S9�	'��a�.���}�݁`�PP1s�B1�q���^s[��`�ω����1�!�6�?bĀ<�3���ú-��)_�Y��G�������M�>����Sz�Z����{Hw�L8b�35T/�R��*ŰF?�r��8��lrp�+�1Q3�tQ^z�e��/����&����rӀ�cp0˪3n�������֋/�?��_��?�岦MC1���*��%.¥OO�ɋ�Nh�Y�����E�=��$&ϩ`d�+�czl�����>^������}y���۽-�������Z13ɋ{�7"��g�A���IA:q���9V0N�Au��Ҩ�Lr��v؄^�E�bnx\.�,���93>#�^}F&���G�i*����f�mH�dZ�陟��<s���;oȻ�����6�cZ`�.��⁯F�]�[��\��<W`�W{M��9iڻ�R�+w>�H���1�U	���/m%���?+�r��8�����0RP��@ۜ��'�5v�vs�]Wm���Κcybb�̐�8	���%1<">���tc���"�ve8��1���n|M^��w���,��w>�-�ޓb��\9Oʄz93�?%�lZ�E��Y�N��������~#�ۯ~.��+���W[e�n9����\S�|�$���KW$>:-m4�[f������pV�c�[��lQld�`���v&����	:�fמy`���9'W�h*��w�	�"�F�v��p��$|`��ʡ'��&bp_�`J��Y�a���e~jZ�q��r��EI�0G�%��1� *4r��drbJ����3��D���嫒���#���o�����,[7��3��r�*(9����5?��]�c�{/�rzXI�nX���O�i'Ƹ�̢�	����|��/l��:�v���Q�D{�!��-�T�_���|��E�y�}M�T�95	��� ѳRK��\)���+JX�$�?_�tI��xE�k�u��2��qs{GV���d�@!j$�����y���bK����D4M�����|�ߒr�#����5�ڼ�Q>½��U�1I��tV�HF�2g�NKv�K*M�*K�My�Z�褸�1*n"_�I=�)}�Kh؋���I(���Ы�z�*���,���Y�~��	m�%��[!��`(�L�g�cNLr0��r�!`�$�a�#s�1͛�4Τ�2���!Ԙ�P����|��W5��.�n#�¤|C��B�o}$}|[�{��nߒ|���ʷ^a����&�U�ƥ5��dE~S�q�9`S�xD���M��h�N�sf��_���LPX�r���Y
�����������l �E�R,���YO�0�A[��S>�D(�]B�tC�������d �GAa[�r��J�54��8����,`�k���=�|���i������V@n����ӎd�FY*bZD����������a:Fe��K2��	&M`��0�r��G����=��G�h\��
�tzq^p�����	�s�����J�_>y]���fEW�j�:��i�*`�Z�䠺��<�����7	���<PE=��7HFdl(#����;m�5"�6h��t��&�H�7	��v�9X4$��������Pե�b����8��/��j}}�7�,+&�am˵J׫_�������F�;�$�4n���t`�?�|���_�C}X	�d����ǒw��y����\�]��{�HZ����Ƥ4�Ώ�#�;�h�%w�
��Jo��l�G��|OH���#6g�0���AZs��_�C��-��<{Π�>%�?����샎�Uhb�.�z4�0��Rפ=��B� �d<.�g?�|��3�Ԁb�F ~X⚟�A��u
T|p�""ZS�y�GdjnFҠ�P%.7j�QY�:�$w�d���]hn�0mGR��g}���<�1��n�>͌�8=�j�m!�	3���;�N����&d*PF�:6���r�Vh�/956�+���B��r�fv�<��\��]M�l׌$�-��4M�Z�W���|#��1K+P'4	[b��'�D]��q������T��\T������MM�*ǠE���dh����=�N�ب��1����}9}F��i���,-.�i��+;[ܔӰ���u�;X|C`��K\�z����^p��)eҨ�ٔO��zA�W� w��A�z����� ���{�s��S���
���hp���S�w�1y�1*���փ���KL�����(��ƸTY]N:Q����&�~x2����Ou�����	���eye�m��]r�G����<vva^�ΨİL!�񾌺a5ȧ�fu�W��2F<�iJ�p���!
���l�w�6	U�"}�	CX$Վ�0$��#G	^��yά
諯�$��+���J�I��z���%�/KC�jQ8�KvkΩb�"�����5*�	�Lq}�հu������'�z�����k�7s\���Ua4yF
����JI��|�?�#}��=)�#�R&�w��Aa)4��979)�Ξ�Oޗ���v��Z��DG���#7��B��f���
VL���Wv�����G�
�gY׾�h/@���D�\> ��
��A�������Q�����?%7�'|���<��<�����kE��n���߄�\�2{H̋]��CC�*���p�#g-;"��?��1#a�yPZc��uPP Ϝ��V��4!���ĉ%R,�aO�����m[�q�9y+�4np�(dOc���yVc�&�ًGj4H���w��9=�G�"���T��B�q;S��^)a�Dν��Bq�Y�eD��������=����H�T�sg��_��_ɝ�����d���U��T�Ǩl�� q7m�U	B�o�Srnj^��}%��+���"/~��կ���y��C��ЯQeP+?;1N"p� ��l]^4�74*ן�F:�'뛜�QO��K/��|��Y���f�dinQ��-�}ݗ|���\��Aa0�f
I���W ^,d��#]m�R�Ǟ���qմk��"*�~�oS�>�{'}�o��}ϼR�Hť"�Q��º�Wu}������T�<��S�v�0��BܨE�|��I w�Cb51y��f��d�����Ĉ+�]#�`��ޏT2#y�ɀ�8E� �.]Д��T@��Ҡ�p	���C���359}���@���T����6�JjJ�=����Ь�|8AL���W��Z��Z9+�6W�,w��WU��*�,b���P+��0�����jC��K� �	�I�y��i3b�H�/��0��iIʖ
,��\\�\��uXˇ�Ȉs��AI�'�M��`F��&$�J����xŪ$G�̹s���c.1>3.�����]9P��$H�v��'��.gD�p��y�v�C��aS1m���g�� �o���@�3MW��8
��,�5�l��<�k�Va�Im;p	�%'�����kw�_&�[�8!�G�#p]��b�Lh��{O�{���h�,š��y_���'j�@[����ch¿�-�@	��2�@Q2�$�o���B�p�]�x�q� u��!!�/Ψ�z@1���T� �H�9N1Ϛ�����qG�Z;�.�*X7���l��$�,����UQ<�y�{xLi���Ѫ[��{�^�@�+���/��y��2��C3�b�yR"̪�ڲ�������q��P�3gN��|�v_�阔|�4i���FmV�r��:ܸ�CS�Bf"B��K�/I}jFk<>41"Ӌ��oT�]�'�T����F�ɵUޘ�������~�O�x�	UC+�������7ޠ����?�a�.h��?v(e_�yT˂ZĻk�a�g�-�X�*�%��|��~�i[�"����V�i�z����1�<�u�,����Y�f8��GQ	�
;SS֛\���<���#��c\����A�؂ϡ��w��8\k�lbY�FZ(�K%X�9��}��\�n��	��w�s����s�5���=��8?t�V�w�;�8� �F%�����dc{C�_Q��N��x:�S���}9^��VG�#���r�� ���Es���BnK��$��������2y�#r�\�dI��$�,Đ�B��9����a|H���N�*�lRb����}�l>�{[F�a���e�`[n=�'k��L�;�7��&��j$��%b#��ck��-������Ώ>ԛ~���˪�/�D�Hx' ��<; ;�!�z�z�aM�[��A3���.f9�l�ZI�@z��*`ynj�Z��^�Fv�������ӯR_�K�z*��>_x>���)	�<�R�7;f���g��z��=��`�$M���k�_C!�S����4d�����yc�z�ww	�+����]6�OiT�5ۘ��1���as����IJ�����=#g!oL���mb�J&N�"�;*J�ؒ���rMC��P^J���Q鉄2Q�f�����^�*�#rP��U+R������.N0� 5Ċ�Y5�1k�R����g%�'��Ȅz��Ȁ��i՚$��p�/%6��. ��;H���0!l8�ĀzA<p���Y�����͏>�S
�#b��nsg�Q]��ަ������krRY�78:�͗���ן�;�0�굫2���W"����z��> L��JebH� �E��PrlNM��5�L�i�1�>(`��JV���+hL{���]1��G&31ś^��vM�}�=�~�\H�����ۥ����G��S:mfRp]�KA}�S<{>P����؉nv�K4LL�k�G�gz�+�y��d�6����E��k����q&��`��t��6��n�]F�������B�Z�J� 1��>s,Ɓ����$w�Y�	_y�e�0=�u��o}������K�^#�u�.X\A[oF	k_�T�kd��,�$�{z2�����	���c�^M9,��	�.�p!��h�t���j�.�olIՍta4��zp�`�Q	���x���͹��e��%O� x�C¶���2�
�N��'B\/2��a�0o�%꙯=/E�`�ޕgn</W�]�S3��[V�sƤP)��a�[i]����ݗ���;���i�U�ivvV�w��Kh��� ���U='���>�������[�v&<�"x�����(�U��K��}![?�O�3�$�}L���������;K� I����Q������v	8O1Kn�@�o�x��;Y�iIbaunY޿�#i�^��}�UY:wV��p_���on�ǟ|"���ؗF�8Ot0u�܍2=5m�<� B7;`jW��v�R8.�����{�X���qR�3|s�@�ܘ?%�յNd���F��S�"Oj9���!w6wd=_�u�U����������:��3R��M,A)U��䤜TkX���چ�z\R�>)c2�$�;-?bU���@�KE-[�ӔɅ9�[���Z)Gs��~-�r䋉9�6 Xn�����iɊ�������$�!�p (���-*��?溬Uz�YX\\d��\W�^�c�� ��eugS�}UU�Nzj����%�_���	N�W��@Ў<������K���D�F����"��pj��h��)G0����`e3���≊�caa�w��?٧Z5���v=N���ژ�����X�W��7e��)�FT�NVZeN��h����FED��ްhk�1��U�N�)�5F��_����,���/���@S����[��wTx�2v����2���� �Z]��-9h9r�@��J�Ĺx��b�A�Z�|��Q+j8�D��߽���4|�<;ϭ��اwS~s��A�v�K���&�S3�|X�V��!)5k���H&��kg/��������V�-���febvFv7�0�B!�ïQ����ʷy�/w����IT4tͤS\���˗YՄ���UV9р���m����E���z��D���P߿u�t�y�	G|<��B՗��d�-���w��O��h�gz�^wX�+�����Jwu�������u�=8�͗Aw�`�1ˎ����
���ٽ����i���զ�DQEX������!3�_j���]G&�e��9��� �"]F� 0�}��-Y���NI�Ҕ$��U���'rom��^�����
�JeM�A���T�GoU�˨��v[$�BU�f'�U�(�0Ј<
,αT�4RUX��	����c5��^������l�?�o�pC����w�}]�U+��U���F)�s+��2�!^A��X���@�Գ��^���gS�SY9==+A�;�Z�*�JNY]�� �2d�	zTh�����I!7�Vyd`�+�ϝ;#�����2"�723`h*|�(��?���Ի���n��?��߈��d�Rh���uh�8%n��m�b�)1�s4�H��HmQqe�߶2J�.�ڳ}I�}�S�{����mӅ�-�|��%��V\�7�`%~����� ��q5PT���S�,�rb`/�)�{޼V��Y>S�BѬ�Fːk�٤���l!��ovb��oI�y~]f�r��]�&����_��S9WD����)C��/�*\/ �B�5�^�V*Jn[��%U5"���d9�+����}0! p�5���b�d�#֋د��~^��Z|,r1�e�q�̅q#�"aq�a!/�ۛr��]��F��U���3c�֜�xe��YШ�JH-UD`���r��Ŧ
�>��`Z�G)�lKMC(�x_�h�j(٩Xb!�/
"}J��k{;D���ϰ�{��}2IϪ����#X9�~�|&h��d�p��_��¾����փ��B��Z�H��`G��/O�xH�g߳[H�,�^��tf�o?��wCͯ�q	�$���{�,�i�F3֝�_�P���*�?4�y-�E�|ɉ{� e���k�J�=�{;���p2a �m��Y�`��H����GrnzN���C��O��CR����ʁq��*W�z�`�0X�k� �u՞�Р<�-�o?xG~{���k��|dӔ�L�����K'őT;&�q|�� Ќ��4�VPa��H$����>p�P)n}i�}B2�n�©32�֬�_��<-PC��K��v���/�=��,��ɫ/?'�bE65��5��֒�z[���ܕ����ƞ�y��+���)�,V5TEߑ�V��7���Ԙ~(�f{ ȉͭ2���Ò�4�%"�3`	� g�6*�[ؓ;�����*,`�9�w��:'�ʴ-��J��0����t-��_�N��̓�E��H��񚯧ʝ���6H=x��F�j�G���S��l�(7m�=�jMl�m�Qߞ�0��`����RRq�҇�i[ 32��2�@��d4�)�'�żD���w� �nߓ��� �����5`k--H_H��|qu�T�OI8��yF~���_�?�|M�*R��vǾ�_��g��ICU�*A��/d���e�{��	��E�}�.bhP,V�[�x������(~麆�9yc���][�'����|	;�;������>'�#ϝ:+G����o��?��PU�U��p�Jd���5��xZ�^�$�g���[�H�P��8��اPՐ%¦�Л��}�(>�/e��W.\�S�Ӳ��#O4��h�`'�� aB(���%/ߖ[���z���e����!�cc�M�D����/����ޤ<O�|}���p���W��}G0�i6G^�+za��J�i��/>��1�R�=eCų�o'�7��@�Z����@��*7��u
q?R T�?j\�<��{+�6<O���$=.�U`WßIӟL��g�%!�����ir~������?xW6�4�>7����N��8���e��F����ՠ��0�iK�e���9��a���?djzR�4�8�ޣ� �r��r���ǋ��o��d�;/}K����n} ���e3���>��
{"-v�%��k_ASX��ե�rzjT��6�����қ�p��LNͰ���=��˗����7?��!H�u��ї�%6Mv����'�oJI�ҥ�%�(�t��]�}5U	S �QE�7��V�kG{��s������C��E�8 v���K����޳X{0��A�o���ʥE���h����a�>]X������c�K؟rz���,�+��%�@A����d���Ή�1F8D�rA2���nލS��&���ȧ[$AN����s�5�JXݴV����xN�b������5�lzz��-I�4�h:|�<�N�!k8a��*��W-�K�` P�Pc�ԜmHS@V �n�[�AC+y�R,.,�=�Ͽ��V��/�HV��2������!k�ǆܼ:z?�R� �O6SY��R�ۆwĠ4<�;ɍ3}%b[�2��	d\bt���C��_��2"`�����&'�e65 �&��Z8%1�h@��nܗ�G�j��>$dq~NΜ�����V�$!��)���
c�\������(x��>,�5���,��f#1�!:�z�U6�B�����-�%W,HI��B")3�v]Kg��g�|��� �tn]�&�h��ӓ��|��u,�Y������|�g�)h��T;�;)�?���$��ʌ�
���&�I7��U�J�(>�~x�`�w�e=/�#f�_jn�L�Ͷu��\�z꿷Ty|xD��,�m�񷊞g�p$#�����*[a)AkE����a=f_|�E2��ۛ����-�c����B&�/���=���#	(J�כ��Pe@ɠV��Z��T��/�aU@yױJ(�	M����^|\�9�����Ʉ��U�c�-N�Y��5�k�Y�Ҡa�O�Z���bj��D�[�0i��}_�O��mdNa���"��a64t���=��$6Ȑim:XB,�(hR�ˑz�,7���;�{�!6�1��#�JHG����kP!�3�}uV!�(����������fx���D0���Υ��z�g}��:Oy>��{���]l��ӝ�8�����(O�ßŭ�`Ja:~��A�^C3�����
�B�2"��
r>�<�M���K>768��w�}Lϒc�h!(�a��a���H%��[R��0���\"�"U~R����o>|����m]����O嫓ԟKb�0��s�Ͻ45aU��^Ը����I����dRѯ�Uj�������c�8.�N�%u{U	FJ�>������nL�ܽwW���W>Q�R/TdxlJ�c��у[�}�O
>�V�U9R�~P�I�V�0�w;2\ËeX\�M���T���CIт��sG��.��/.��zw��m���Vk,�sw�R��Q�q|�%V^�bF0�d��CC����*���L�k	� �dI����Q=ߐ�Ah�b(����� �{2��*�ӽ֓�9,�
��G��#�&�Oz�$��`��l��
G����g�������A�>�3�,���W��[��
���\��C	<�{&�l��;fj�7����%��(��P�q�9��傴5E���YHD��#BLD@P�N,bWʙ�%O0L�n���E����߾�0#�k2�r$�hCB���'J8�
���#G���vrK�ɲ����Y �C�$�sB�ñ��lk~����?K�H�*�,s�����:���5����G�{pI�^Wb7"}V����t���8  vi@w��g�+IK�W�h�<\i%`ER��  f 0c03=��+_�U�mD����/2��z�1'��dEF|�=�}����'Pi�uf�f��Xԩ��$j��[�4�J�)�2�]���c�pek�F��O�n�>u>TwO]iGE���/ Z*J�J55�� .Sp+�N�c#@߿��o��s�T8Z|��Z��@km��C-�t:ŀf\�<M�$�& .9��XK�X�o���C�z\���&��=��Y��{��p*FzC�1�>q�G��+�`pa�'��Ece� ��O/�f�ō��|<>��$�ɱ�H vwRb��g�6���0�����i&]��c�C�,��=��C�z�Ð�LYi�Mg�z�O��}f��Qv����E6�@���)yп��'�?<�k�]����nc6���`��s�U���&2s�J����nk�MXQ���T�� X�#��?}�w��A���+d���v���qq���ؽ��gN_P}M{��*vE�I̢7�sY�͒�r����o�;Gp��㧌�>C�V�/9{�I�P1WT�`��V���	�o�!&S�Pϴ<�je����̷�x{��K����@���͒D�=�#đY�(�
�1����
+z�;�M������p����G7�����|��'F����_R�4�sȝѽ�Ȟz
xH�T�S�Xv���N����>�'�ɞ�`Q<�@�I=2R/>3.$6I�z����>P�39G�?t�����ħ�yb
3�|��x�~�R�=���'��r�k��~.cf�N\|S+KJ���[���%���8;/���iT�
��������3�4�i�u8�ab��j��t�^��"$�f�B�� `������֖��SZU�-ZAm�E�&�]��6�ެܛh�A���M����s��{��t�(�Ʌm��s1c3�����̃s]缱_��%.M��;2�]�`�����R�3��_f��N�#�(���Q$�m��{8-�d3ֻ�@LZ"�`2���FTL�կ}瀏	}-/�3�����59' �������=�O/}�>�`��y�K���Cw�&1��X;q��@���Y]���º��c7
|4s^�&0������w�I�ab}����Pݤ�/���e�e|`��;q��-l\���K��'����G��n����Oc��1t�����h����	4&��}9��n���ݻh�#��������qR��E]���>g;����{e�ժ|��g�E�YjX�H̲�頖���@\�5�y��GS+�������AW������ߝ�LZ�y�l�&8,y����c)*�=��`&�	��b�)�ł�9["x��ZyZ_ƪL&N�L�KL���L	��#p��t���H�� 8���߬��:�-c>��Uهcn��P�N����[��ͳ�7c����Cd�6�a�]:!9�H�'�;��f-�~\��!k苙8���g0p#ͽO�O���p�u���:q�`�u���^�'����
���Sg.��ӿ���:����97 ���T����R�خ����n?��[��E��k����Bnx,jg�y��_Xė�x�fgŚֱ�S�͍Ul5vuߩ�'0�+������|�����Ja�h�9K@n�EӐ�3-�}u�W��"Z�~�����[���������s����{�7_���	�w��ӷ^�߿�����L"7towW'���@0S��G^K��Y˼B�d��2��D�Wr����r;u��-�E ���|~��wF@��@����YSS��N#�vu�w6 ōK���A�8�A[$��A$�Eb���p�$�Z甗~j|�Sa�f�����U�k��Sh&5�t�ߣ��zK�rg$c�\���a[]�V��+��:��=��$Җ}�s�z��X�a��~�(�N}��	Q�9L͖��)k�!>����<Ƒ=Σ��D�d�{�L�6�n���&L���Bz6������ژf��!�"S�
�Pܟr�S�id�e��6q�܃����E��!Z�mҔ=և�Q^8���X�D��2F��Q�:�%��un`�\BjD"H����xT,n^6_���wo�/>��������ߎ�&/�����)7�ϕ�u�D`BN|�'�΃����e*�q����"�=}��e#`��/<��f�����+�M��E��n��'0h��C�Hδ�6�B���y7
K�u�9��Ğ�a
�9��o���{�8K7��Nv�л���U���ϋ�&Z���ݽt���9HE8��jB�6��2�����ί�f�ϗ��w����������Y�H����~�c+�+��^�jv���
��a���_��Wp���n�h���"�l���v�����۬:My�ē��.1n6�.F����\g��Z��M!d����m	��$ ]	dQj}L�gP�Z���h�,��>�wY?L6u~Z�Ȓ"bY�R1�ɉ��U6T����lC2�F|�Ti�2��2JbYI��۩��^���$NN����W1W��<M�����ѩ���ˆƝHW)0�[7nZ'?;c�?��E �y�#6��ZuJn�Soak{�Z;b��)���G��ͫx��'�a�� >�M�����-��.���3be	�!9x��f�8��\0;;����Z뛴tr����项��lhW�r��N��A��JZ�k�Iڕz>��<���BLW���zQpH3|����,	$.#�>B�x����|�P418bԳu$rIg���Jw��:r�lll8R偮I!���΍m�Z���^�ٵSx�G��铊��3��y��b����U�g%�Y�ߜ,aG�خ�%���3��2F�x����.���$�˧
k����	��ʆ��%��lys�Y �����R����aqP��m�a���M��_Zͥ���3:�=yo@���o��&�����w�_F}ҲgeC�.�������}AջS�bQ}�Q\x袢VVVp����q��jڋGQz�_(�ғ�<���Qa>y�B�.��ݹ~�~G,��2��qA���蟼�fZVi��5zH��X.`�K1Ʋ��{�Ř��"�\LB0����UW�/q�0�Y��W�I6kj�"�D�u����DK��4?�M
R��h��a���3��tM��}�ә��*��ص�l�Z�Awn��r舠qH��֦2�g\{-���}����Ʈ��l��3
��z���6E� ��\b��������'O����S��B�.agk�}l��^v�������Y��sε��M�p������h�@6ms����!~t����� ���}#�������qB�n���CQ{\��h@��Uk{x�o�\��?}o��&.߹��N�TIk#E��	Ĺ yQe�4����#:�O�㖶R6��T�෾������%����)�tS���Q����_������Ekh�%�v�Ct�-Ea����x��7P�:�O��2�k��p^!]��~I����T�v(f�8Z��5KŢ�&I�Dgz�Z�"�21YHɄ�зԌ�6t3m]���|@�䴘�-�b1W��[�5�M�/%�I�ȭ��ߌ�9��c�e���Nг�l{��5Mι�с��+�����y�ϯRW�*RF��d������;x�g?�믿�ύ�C���7B��:�ͱ��}���Z��&���ng`�*�=��ހ��t�]�.�2v�qyu��%L�>}X��g�a:���v�Y�&C\��[� 70^�H�+QyQ�W����Z��.
�_�n��VYϝn��9m��j��&]�6�T�����������E��k�M���L�i�	_[�o#�k� �q;$�͗%Ԝ���&�r����J&�U���@��{f�]d�@�ekoO~�C�t�x�S3�s,�9��xG��k��7^C"�~�X�����$NN?��fe\�qCq���eq���K��Ӥ��ٗx/�Y�9�ʭ��{�q�k�`A�����6G�%�1j�Ai�|�k&N���Tvm���ھn�j�@�ljEO��xQ�2�+i�\q�.<�B����L6�z��+�v��rٴ����I�9l�"]���6._��=���EM�4��v�f�x�����jhB>���l�\�<+�V&#+��~�ʫ+�we��D�v8uY��SgO����5,_<+{��w߾lJ5\���P��n�%��m-�8�-&�M]��q���ǧʘ���{����d��浤�y��	���{.n�˵�����-T�J�].�g�����2��)_3ӧ�0�<�g�e,cen�n]�~��R<�	=��֏z�/���&��_���K�-O4�R�c����vs������呫�Ŧ\��D����%��� �m��N�0/�@�j��h��i��9�{b���cfm���\�A4�u�`ӏ'�U�"p�ʮ���
������XC
���p��K�%������],�,�nv�t���_�/Q�{)I7%I�_���
�����a�N]ϬQp�#��g�y7n^�����ЉC��.�)�h167SلNI�@�籱;�Fe� oI�ĕ�����?��:S9��m#���~������X�X�Q�Ϝ>��vW�l #q`��u#�����f�O{�Y��M�%1g�Z�����թ�X��Q�{��L�O\x���~u�	[_�Qۓ�w��rs�և��^�v�H{�\�Q��d#�.�g�cf�Z;H8�Dwi����R�ss��4�!��s�ԴhS�3�H��ٌ/��>�������sX߭�h�&�׉4����&#�3u	(/E�la_6-)�{e���)�t����X;qM��T��Q���`���FQR���$����#k�Q���������8�~>>Q���'\����{?�`nvN\ʲs?�?�V�7}UJ6�y>���z�Kz����t����yb�N��m?���^Ӗ�vw�����K''yNN/T<�f �C��������P<T�tS����8@�4���,J��aV���ݝ]䯊w����r��r+S�����1�2��2��.+7"�
��l2O�R�)�F�@7�m�_[��S��cE�Yo�6��w�"�=�0&��N�1ܽ�����$[5'����V�;;Ml�˧�J�,�n�ǉ���1HA8����Z�P~�J\�<�k��*����(x�C�DX�󷾅?������[Єh�ɹY��wwdQ%v�k��j/l�HO}O�FA�xGY�`l�QуFe�r���,f�Ce��6�#�b?' �������;؝O�k�֭�&>T 3��š"#J��Ss��T�-N�7^7{�H�Ө75�ϹdF�>C7�fnC���5cݍ�f��ks�iaY�W�Y[ϐ�7�'9|���I�e��u�+tN�<�p�!�T���!�"�.x��p����9~�����H�EQ*P;/�������ZSԽhu=u<X��b��a�/���+c�`����R�^�Z�6��F���E�Xr�V4ȧ�?;�HJ��r���d#���*�0���%vh��}��� `KD)'��b n_}G���Z!^�Q��nְC�a�~0Bv��L2���~(��"%��<t��հ#�D��._* Ͽ�Q#á0X�J���\=���r�&����e�C��$�e����ډ�Ќ���DJw�P#�G$�9c$N0�^2D��n`8H�t,.-���P�����Jŀ�y���5sY���V�WBZ>0Z���#��s|#E.��KEaa�������_7�B1�3�#�]F�BA�ǒC��SR�_5���X�3�q䑱f��wGc�g��{NUb7�(5�9R��N��\�v���0�%v�n�����!\7�>��V���m��׬uE��K���J�Cg��ie�u�;BC¸�){���DE�WE^���ʅ,-��ˑ�1�7�NQwMY�=qV�^���Wo�a��C���$�>49���̀�� ����2hCF�D$�����͔P����J�����`��=�*r���]B�8�H:|Q*D)Pp�8�&���,���������·W����;�m��Xt���Ąā��
�-�A.8b�A^�xܬ��uc�r�=���ǧ�39�6�V��"24�X�X��ۍo�C\_vL3�ݭnk����Q8�6�W�1���79���<#J��h��9�Ա�������Wܛ��%�9��{d��P��&��h�)x��IG.�6��u�u�W���� ��F��-�˞�9{���qbe��4P��4kD����srF�W�q���4F��h��E���hV�����ϝ8�S"���y��I[�M|pgW���^`-�b[6N_A���k"M�l�-���8�R��ڲ�ج;�){�.�<�����0�������:S6Dh���E��(�5ȥ���:�NԔ��f4(,������Ν���=����ΐ(�.������3��&���!��'���D�5����ҋ�cB�)�u҇���Kx�a	c?J��m)�5��ڌ(�"(�h�R�	�o�5d�Y��e�����M���ɹ��'����̗ ~��Z�\�C�x���.�R�wV���$��X<�p,?���Ժ�{���(�����w����ц�������|Y�oQޛ�0+��8�z��V���U�>�Ÿ��B�Ԭ��w'����iߗ��Js��7� �le�"*F����z�V�����ؐȤEbs2��2t�5=��m쥫�6�{ea�������|ss���֝��Y[8)��Sg�y{�w���]mU�8+�\')g�!TTk<��g��K7������rA�b�z��(�C���}���ε���Z���J�����V{��>��A��`I�^o�\"��4T0���� B2Қ����T���]�����!77�k�Y 킍:f-���L��Ff9��(��i���.�dm0�$�˧�����"�䋁���ԗp�d2�y�1��l�k��)4Z�b-�Ą��/���i��DɁ>B
��^��|����_��z2��]Q>����ٜ���J����*�Zܚ�T���X���B�5]����⴬yE�aRG��ױ�=f֓8����#��������<���ʱROX��aU�d�����;�i�(݈���%��>{�Zf�q�{B+�[�I�.�מ�"�����%������70�Ty?ƌXڇΜõ_�������:vؒ��-g-$��$�$�eZC����%uL�Z�:+�w�s(Ξ�I������hȢ��xJ�^�#}�Ջ�v�~|�cH�Q3���7I-H�gw�V?��r^�<d"�\&:�MK�9)l<��Mn *��!�]�0��~#R#��=?F{tܿ����%��w���yN�_���U���z��
f�4
�bGZ�CY[�}�W�R��<S6S��|�B�2��)�E�ڨ����������'��o��o��o[���&�TX7�e~K�J�.�o�e�]�5"�:#�04�U�X�\�p���̸e�M	���ęH��c��v�)ځ��o[ɔ?j&
�2m�i�1_A&^�C+B�|���y��$Q!,�%���U��"C�X^�qy�zq��<��h����u�f�8Č�4�uK�'����^�,aE3
��ƅKA"B׶���w�Ôh�Gϝ�!+5��#c�dY�Џ'M<���]�Cff2!����aU�|R����� ��t�sBm�	aBj�}�(Cͽ������W�*1�g!o�9ّ9��=3)J)�����Q��=��T��:.l?(65�d4�|�ge��Ώ�^;��_���p��i��?��/��£s!dmɨǚ,6�Ø��U��Cbd&�8�'|�<"ψϘ4�|�� �~S��+�Z����=W:J�?��p�@%�!��+YR���X��]>䂸}䟌�o���WJ]���Y�X���pv5��|����FkC0�^��
��]-=LNL���]O`	��qư4�n����<g�aKH��'WJ`�_���myϻ�5kJ;�mT�-���%J�D��`��|"�-&5+k�0�^��`�q��⢎;s�4{�Q!m��y>�g�N�쟾�3\z�=}Ȍe�u�i�]FkDw����/�'�h��Y��w.F;��I6��4m:+��3���}�q�gڔ뾲��h�G�yx�%���c�u;u��|�1}BT|�owW�%��W�*���s�mT���N�w�p6R��l�:�c�j�t�Y��H����r~��
��aʣF�'��P����j~��l@����!2������b�H�iޱŤ�'u(.e{O6��-�f�#?]A�����Jb����������[���}�����HK���ɦ�uZ쉵�!y_+r�����K��ݬqĴ�*nu�p����^Z�u֧ǵ��i0F�Ƈ��|]Ѳ��͊E�{��&y�aT�g#�����أ���÷��m��ʫ6�X⺎l�b��c�ǰ,10�^���_b��Ȏp��x���m��`t�0/'}�c�J_����͵�LL����b/L��:���]T>C��*'�_��r�C2!�J-Ŵ�kt�6j�5�w��-���﫠�g�J�V�q��|�k_exҬ}de�(Z]O���b�����*���
���wu����"����h�(͈�G�~G����'����$���	m�c�O��!~����c`CB����7�;|����e���������y\}���j\�q;[�8sj	O=�8�f�P���+/��[wW�� Ф�X^��&6�.tEl�0�I�����N�_��s{��-8�#KY��?�y�O�G8w�$^�u|��Ç7��C�ã��w0��I�f#9j�sڧg,ڀKj�g�yF-�����ȃ u�ܡ���$����1�����a���s��`IH��W���U2���Fq��m��_�C�/��R0 �ōj��|ĂK����9���Z>;
.�����ۮ�ĕo�E�8�?!t��'��u>���8CY3H@
��H�\�����ydEe=�{n/34���g6vM�4Z`5>�&5�mln7q�u�Ӡ�M���Υ-���_GF,oY��3��6ʴr�QU3�р��y9=3N��*��]{�z�f��]�<���~�o�;<w�AT�"���<�;���o�o]�E���GxB� ��
t(rs,r�l�9(�O=��>DB�&N�B�׍���kh@c&��(.܀�����}��`7�Zq�ѯ��w�0��E����S�H��&�QbY?:Ϳ��:����Nu���ߊ�=^�^�S��=1�̢�[	�~M/�*O�G�~��5\&qCO�-H�#z!�̱�ʭh��.��6�ŷz�}ֹ�����N��غ{�(�z�
e��>hb@H����ʅ�z_�2&��li̖�m���Bq�t}�A:�|�Zx���u,1jN��Њ�<�}s��s?�@��7~�"�[ё�{�W���5nfY�K��U�R����.�5U��y����i��4�ɎҌF*i�_�t�H���\*���/	����G�{�2V�?���f��>����1��>ܽ�>�8���z�T�#���ׯ�f���l�ݻk�Җ=z\����)�7���\oo�a�j��M;6)*U"�#RJ�Q	%�G�2E��B�zE�E�E��M ��V���8�8�ݹ��.�݌��sw7��9�b��qi~� ��E.͟w����P��R�����(�ʥw.)�5�4��S!�ߺ�nd�C�猺�2���n��X#���5�\���y�9	������R2٭_��/}	��ru4I-�W�v��p�}d����r�"m�?N<2�Y+��E��m���S)U��'Y5]�P��'�<�c��\&�1�Y!���H/.��=��H!��G��s�p&v�W��-����bG����3
!3uy�u#�m����>��B-�D������XqޕH�c:̰��\�V�m�z�����I�P�YY��FYV��CE QݚW�ح����j5��e�rBp�"V�<E]�»�G�5Ӻ�0�#qN%��N���I<9;����EИ)��M�4��G�����R9��[�i�Zp����4��� 4I�Pp�K	�e�g��b�(3���K�Z�P�X"5���8ӝ��JO�����O��:w�|�~��K��ڒ�y�t�����ӗ�7_{�?w_�Y����ᇗ��m���'����4k{q��z��Y
 Vt�<���rpp�M�q]���䡇q@<#�2�޵�Y(_�m��"H��7���>��}����RJ�Ù��h��?��9�����G[���Wz�9���-��Q���x3��[���\XX���c|3~Zg}�-�A��r��\'C���.�s��d\M2f�C�`l^�ؽؚ��c��$]	�Ef��~���sOc������c6;�\�,V�(Z�t��b��ʩ9<�Ps7��z�[!v%l)h�Q2ْ�JL#֭����>kpbi��L�B����nSNT��]�K���Qo�릞�c`|NS����,�;zA,��}B�+��2�/<�����[޿q�����ͻZW�O������	�����v{��Y�bﷆGP`���x�LOV�]���
"ݖ��s��t�d>�L>�u�1������U~ⱗKD8|Q���jo��֪�Y�C�W�H/�]K._p�D���k;�:����
u��3��e�(g$�l�^^YNۮ�8c�L6L)Ӗ���}���}2iC/�(��ҿ+�Ĭ'���15��<tw8m����ܤf��h��N�ğ<�,��u���@9*"�z��c(N/�����ƺ
��T����6n����H�gE�hTaZ�%�����o��a.���ٝ�h�F��58P�4���P�����O)����ױ-Z�ښ��tO��~�w����l+f���$M%$�X�)qE�Hg"emc�?�a�!aM�(��.]qmÉ�u�ER�19���V�ԟWș�$�V%��N�Ώ;��I�˅
DПiq:3r;SW*������f�s�%���K�_���[m*QQ�	��)�{[��=������0�es��e{<"$k�ENF�O5�HY�ل.>��[_[O,�b� ��X2cF�e!�!È�ɀ�|6x7�m�C�k��=W���Φn��i���g�[�=��r�7.�E�����}�g���gJR�
����Ѹ{	͍p�8�78�|�!��G����В/�~�r�.��sg�,7p�	t�[9���t'O�R�gW�E^8�?(��d^z��_���A�T�� m�٘+.k��.��c�� a+N	Sb�
�H�В{)�-�>�Dd��v%�k#�g4�	�A�t���fY��Y�8L]\�[�nbJ�qa~6$�(���@��11�Q�{��4G�R$�d�E]�h���I��v�
g�~A��`6�1_O'=9PvtP�
��Y������Иެ�86��Ȁ��B끱~>te{Cu,炂���⇱B7�SS����-/S+k�"��Z-ښ��/?���#Ѧe޻>�l&_D)h4�,W̹�c�U��X�U�b�y2ymM��։Pt��A��s˧�`e;o�'�i�}��1w�Q%ɅB�9��Ϝ��DY6WA,�벲{xriwZ\n���.�/��B�Mt�u8�h��0B�h3�=��SJ���ko�Û�
�
kE,�ɕcjUH�����V2��ڷ9w<�4;��Ml�Ch��'.	c�=N�m��n��	\,��qӷ{�B�d]��
�7��ֱ'��-��r��5�p>D1�1$-����9e$c/��e���(K�K��ȸ�=�:�"&�c��
7M_>�B�.�j:݁���L����Yq���`H�o�� ]��(A
�Ƕ�I�A��M���Ĕ�ϯ]z-7����w���wI%?����e�fr���bR݌�%9��A�s`Q}�6i]q�}Ng5�h(���Ta��;����Z7#�i�-�����w'�Ntq48H�(ΟB��%BPł���K�l�om6ƴ1���ȹ�K**s��P�^����)��=�n]��u$��+�f����Bsw?u��A}ڹ&n��K�:?���.޺�N�9�G?�$���˵2�3��t��kV\i8-M�r ����c؋��w�EH0w��aL�<��#
-ۥ��D�O�g*�td���qO�?�dRLbF5��"����L���KǿUд�'FnR��3s��4������Θky�8���?�qt0Jy�Nao��Y@g7�򘝙Ŋx::'=���q:Q^!}G���=�uj�P�e/�,�N�V��jd��Š��p�iq�)ެ�4i���[�%,&t��u�^efQ$��k�+3�%"]���W0�~U,O���B�2}Whw�-����Z�\�n�:P�^<�oom�!#7��s~>��NM���\.���K�Kuwg��?������juuo*eL�7��}�{�Xh��C>ozq�r���v���Qd��Ԥħ1��aD�[��]g�[�&�%�/j̚�ӹ�}����.n�[�Ed������$C7H��mU\e�V�{���޶���H��p���ǚxCuӽnK��kc�H��������{˧벚�*Xah,{i΢�{*CP���ژ�2�B=?��|�=�L�Z�#=����礆�������*9�>����,1� %ѝmmF�5�,v��#Ia]]���A�f�B��p�j���,,0�����"����ņHҁ$���0f1�b�e�\�@���VY�6r|��I9[He����Z'$ɭ\�fmA3T�|M;�?����������+�D���������~o]�P!c-Q2��	Fi�qh�#��X2��������`����Hcl:4�7i#)��$vE�%q\��I%��Tp���y@i����ލ�\�_�<������9#Q;Q\G�/s���}�Pk}�&� ,Ӥ�R�m��u���{t�D��$	m����y-'��D���^S�b>�λ��܉S6�WTs!4�a�gMljl��zc�k�nޡ݌�14�ﲷ�n>}(Ck��&�o60��bP���kb���aO�D��x%M�9"Q�I��ٮ1^�Q���w��c�} ��4�ƣ3����eCJHP*n�g��Yy69Vad�Ov#��i'17��"W,�%�h��\�S(J캿����lll+q�apr��1N�p`*<9"��=k��ė�������gw����6�G�s��u53�u�|0c����Ǹ��Y�oԻfm�F"��})�,�=>ɵ�k�kl���� ��"�yh�N���뭃�C74��W��Z��0P�_=��^�_z����2t��1�UV�2�^�j#p�IZ5��P�{�Ӭb�{��w��6��9'���
,��0q5�v]7H�dŪEh���7pô-y�u��Yb�iO����gD(k��}m|[fzB-yX8����(]��HJ� M4%n6JƲS�`FT�������l�qgu���������޾��RH�%2���"+Lɨ�u��:h�f.��9�E����P3�+��x^kG�Y���v鳍}����A)��n	"�@�m&�����I�0�a���p�2�z䀦�%c��!�κ�M��S}���̌�-3t����6�8�3�L.�����8n��8���vxx��t��b>>,N�bO.�N���g�P���������q�|���a����pcu�t�Я�ꨦ��c�����:mY�!8�<1���6�ⶏ=s-���@Y�Y�ڽ����zۉ��	o��Ej���l�3���1�^���~�_�k?���f���B����Yfs$p��q������d|�2���d��ݓ+��w�&b��hp0�L&��u�1f�΄I�|�vv�u�gQ��t����w�]��R�o�Ѻ$8:�sD��0�f�/�������@�	q��%[�yS���if�u���'ו��Z^�[yX Sn'e�o�!�EY|����5�lgq>SARo�֫?�={�7 �h���Ǔ����Bg�4vo�����.��D�|$Q��MA�k� ��F�7P�O���|�L�`���A�\viB�z�nOg�e���v���B���}d�kBAdG6��J���'k��~?z�U�twq��I�w�pW\�v2@�c��űQ��s�W��z�V�1�$�҂2���}�V� ��D� ��r��J��2^#�ruY{vLg�n0��������L��uҮߑ������:�n�L��笸���b�����τ\8j���u<m�)��>+t��P�mI��a��;��u�<95���W���("
H�Q�{fY�ϓ���@���3g���H余#2Ƕ�;�y*�Ϧ�K�Jj�ρX#t.�w]�9�(&���(�|�T"2��^��tB�ϧ�'0�,/������Y<!Z�2-~��ko�D�5�}�Y�����DHk���m���� ��b��hl$\���S$��cs���ߣ{I��&�Y�i���5�߳�'��!9gd�B�p��>��M�aw9����.�?�řY�ݼ�^����栏]b��bw}C�O p}G�ST2#�é'�}r�*}D��=�Zt˴"�D*>jO�.�(�5�й}Y�{&x��g�B���<Z�a4~ɇm��bJ%����)��󬋹?R6��M{*�Z��ߑ
�/�Y����~g&gF��1�aj��i�p��3iÒ_�T��sy���W^��S�`�L�
�#i6�Y� Z*MJE.�wX��Θܳ)��>�3C�,��F��3q.A?��V�'f��r���������}�?�P�����e�4[��kl���$?�W�������f��¨�x��^�j�d���K,%��cc�����{M��ʮ�8[EP�bisْM��,��`���+���u��KE<u���w~%Y����?�{��/b�bz�DO�1��$�*a�#���C�Ҽ��؝����FsC�����.�=�}˺A�}�{F�]=�ùbxơ4|=s�p�ũ��54:��>{�j�~D�4㏜��o���尐y������i�o��[e/�k�Bܵ֫mPLE����rVu���`�s�=F�/����s��*�B�ș��_�M2��2H�uH�G}d�mc�
Y��h�N���Q<#&U4��t������L���P64���	lu#���x�� ����)��wX����>�	���Q��(�Y��+�:%֡ �'�������?��?Dus����b=�|�all��w��wh{�8y��'�(���8{�4����%�N�����m�]rX8��咾�w���j������q�㷴nĀ�6�!�#f��hvZ�S'O�k}��Hc�5N��V�L�p�k��;ʦ#��[��Y����M}�����5;���R�hi����Ļʇb/u�ц=��u�G�Pk�?�Q0w��:����AW��ptǮ��3�˭�7��{����;y���1���"�Ʉ�gF��=գ��pvH&�&a�oG���6����6��&R�+�������Pųǖ���,2��g*"��QF�Y۲�~���Vk��K���P�f]�[>g&�}��'�C�� `<3�̼��t�&N'�����SXW��/�K�<��3�h�B�|.Q��Ib3E��W��������������8}�4>����`�:n�o�0;���֪A�P5^W\�.z��Q��a��Q�fH,%�;/
�p6>�؃v����G?���q��I}�t����~��U��	¨�8�O0Z̵�M�j�Q��uT��M��yH0��+��YY�z�/�m�8q-��f����ާq�+R�8�R���p�c����(p��b�����>�1�Dp���0�{%���g��Vt��%@
b[��ƀ-ڷ�P�4\TtKu����=�N��U�SnС�kr�N����H���+��;գ�	]K��Z\�B��|v'��פ�ocpk��'Ye8�I4#�C+
q��B����~o�&[�������"{�1L�ǭ�*^�j�j��ׅv�+Ѭ�Ki]���G>_p%a*S?ح����1��zE�G"X�����<�S��:e��7���+l�EF��cs�=}KsؗMδzs���1�,p�VS�gc���$㸒Mb�2qDQ1ܽ ��ÁQ���i�m(׮]��Ζ���}��	��,kV�	��ke3E�˃�q�\��K����[U�b-���)���8�?��t_��?��?�x��������fB���]�����ޓ�C���)�J֦����n�ā���Q%��O^ć|�g�yZɮ�FR)E�r�����%<����Y���G�����bƹ�~
�g�t���� �=;�&��GAy����Dr�l���USꆂ�� '�ɷ1{iG��!j�>�D��g����C-س0�1�=E�7���)�`��"}��䬩�$����s2�ڰ������je1����~	�8ѹ|��"�rAN6i�4�m�Y�~=�xC�3�4�b�����R%fj��?�����|�nׯ\ǀ���he��0/fI��O�<�A��o���|��[7���}O�Y���ٸ����8v�Z�[���^�l��>��)�H���T�[�H|�n�x��W��?ip�R�q�wP�u��>�>��K��7�������"�ddW �4��w��O6���uU\��.�~�����Y�e$s#ߘ���Ћ`u��U�Uk�]�0�j��W�q�;'� ۾�<Cs;mě�0�3	S����׻��N\C�L8뛄�1���,�}v�:���6'uu��0�����qT�x����p=~�$�H��4E&0�]�u��ϒ��E\�!�Ht3�:��&ͅ����� ��}ܒE+naf����]�w`�i"h�q7����!��Nhybjf�ˋ(OOj-�Ŀ���(z̜��>c�.��D��j��Kw�%rp2�E�d�n��:j�83�#Q|P�����ݽ����%�6�/�K->Ř{qQg�S[���h��i\"��S|�P�"	Lb}���|�Cb�ꦙ����/b���O��|�c-Kq}�1�f5��Ѿš���5Y���n)�mƑ��F^�=q�=,�e����Z��{=�s�!w`N���c��YU�;���[[����X�\I��-(w�Ƙn�����_�H�!�Z�U��'�i}QY����#�����u$-�\�v��B�舲\|��A����Ιyq��#���G�q��)�  ��IDAT�����B�d�̡�K�zc,��h�d��~������be�ƻq����$��85֖zWus�^:�G�^�?�ׯ_�wn�������촻�PvnhRϳО��'�y�P�x�QK��py���"�������7����)�R1�ٻQ#,Y���]s,Йy7W}oo�`_0 9ݥ�#m�&f��v%�8�֫�!c>jʐ�0GJ��Oi�|���i�j{ޝ�H�SP�x�{����|���`{Ҩ�;�w	#_���d��DKi�'19����4���m�������):m�5�q&��E�\3�}���S'f4ΪUO���bV��dYK�,f��N*(�9�y��?To���a&��ń8�IF�H��q��o�0��ơ��𬈚(�+�_)�TXh�rE�oK �_Gee�z��&�������#�1��G�B޿}��_���F��=��8��c"�UZ�K��L��buo��^�|	{��J	��Z4ŚWEsFva��Y�|q����u=��L���"��� ��C����Cb��xH�>ug(T�ۃ�Ɯ��k���u�Ζ{�F��#����l�~�L�c�P�&
'�#A־n�q��4;:�)u�wi��n�L����ýP5LRԤ s�}���������#�<����)&E�������߬f3����6c펮QF3�b%��u���H6�F[zqڀ�^s3{˧��� r���a,o�7�������.��<}Ԯb�2��eM��3��<��a���zm�G�vq��cGZ���&���]�8&�fa)x6Z9��N����D��&:⢶��F� �%n���©Et�=���^E�C4�D,�����"v�d=R��&��u�;!7.��GߚX&
�f�.��J{A��7��o��ߐ��8���q���n�!�;�3?�C���e�	7���kʍ��#>����L�ϒ�	6�z^��8��S�u�4�v?��1��A8���F%y�Q��c�_Ǥ�n������?�s�P��R�s�q<N���,�'n. �ns�38�7F?j�^����ӌwO�m�%��XB�AV�Pk������N�x,�]D�iW_|������~�6+�-4��D��N�g�h���|sc��1ΜӾ1�����l-��,����?�$����8`� �u�{�DA��aR`6{�n���M�I <UP�U$�����7�6�.�c�p6���cb���2tH����=�����j��h��q��%��̞��,�I��ZW3̥|!	˹�Y'|�Ϗ֑L��I����?�]��{z������M7��O41QQ�S�	cmƾ�x&�홑 �^�qb�Ƃ�`����7@W��AGY5��%�Geǹ�]Ml]c�\=>.)��GdH%mY��uM�TB�|����(hp�h����=���AZj�O��ZoʕC��X��l�RV]䉾�g�<�>F1�ii92̀�p�m1g&��nkb$�F�z��$Ho&)d��C;�{(H [fSnD�|Fц���E(�� 5������Ytm�5�<S7WH[��F���&��W�*���O�;����e��;ν�X���9>�uʈ�8dvw2+�A69]Ypn^Ώ 0�|��?�e����3�Y���I_���f��%?��C�tc�u�X���5e��p��Z%W���$:�yb��LR�ÃQ�r;BZƦ�ھ�t�q��1бo�I��#�Y�Z?�O��{��W�'����$�mS�kW��<�x�p�xa��YRuS9OP�x�����gK�u�k=<��5YƔ��k�g��2�����T�˳���DaU{	���Rk2��1M~x�����e�an�1�*/U�l�EQ�Z�:�8��Ξ����hs0��6�����^����a &�z�z�����i�8m�g�ŋ��B��Y���󡢍���-LW&�<5���C#ꣾ����d�f����h	�F*��)��.MϢ9������^�3s*̫;Uu��0:��ؼ��� ��D��F���0w7Pm�J�q�%]���&�l:��oW_���.�p �Ӧ�	���4I2�������_\��c�g3�i�&�SSX\X��Ң
��}�͂�{�����^�7��er��������c#��:�QqW�@r��;��"�ʚ�sm�6�\���W��-���6�ϻ���	���[�ƅ�[F�t!�R�IT�"N[��1��I��B]�������x0(���4ni-��>?�
Sc+�g
��������>�'g�Q�U��6lV傆��0����sm/������ꅨơZ&�m��9�\]G�D����еd.mV��c���J��|ӓ�XY\Dsg��@]T��M��A�hY>�)�����
�����"�-õ�ۨu�A��1�:�/!���	3a���"�s�ID�<__���
�#a�����k���t�h���P&N�Np�����:�=�^���3�}�k(���+w k
�v��Z-i�B.,.h�_�f������z����7�Y?K-q��:���6=ۨ&p��<�����⵰vʘt������xwG⾞�q_��R+��4����~N�$!�\=ڭ.��/��8��&����v�P��i[�-��>={}~��*��	��{L7����ۈe�-�����<�3��W��+R�M���<-9�j�г'V0!6�|yU~�A�c��}��\ഺfݦX q#���O�F3�ٖ�Z�8����5�|��lW1���s\D�b/����[���
��x��x�?T7oRbH�P���[|lb�x�x�x��Wp��M<}�"����c��-|�/����x����7~/��s��?��s�O�H�"\�V_�>N��K�X"�݄�{ⲵD��jwZݔ���øQ���ؖ����� �?�nJ�yrrJܳ)#Ft�Ȑ��q^�w��Ӌ�g<> ��Y�|�����i�XlccC� ��_2!�!t�L�V+N���Y6u5csz�g9*c�<��X��J��-L�Ģ'�z'�,���������Ɠ�W7�Z�)�ү�j��.ymU
RA��Z*Ϲ��*�,>��:�d7�7N?��呋8��swW����Ϡ2�$�Y$1޶D��"�5��+a�K�qa��>Xå� krd��E\۽�L��)���l��}ufy_~�q��s/u%�[�©����}ӹ�&5��;�����_�
r]eq;����K_����	���;�y�|��g�_��޺���Lv|����|���H�(fK����K�Ji�[��z�״j�Ѳ���"e5z"U���y,+$NS�RQM�~���k�.Zz �Y���Q�p�x��S�sI5��X��μ��F��oV�s�fgtDq��N%mEb�ojjZ��xS�=>�tp��O��=a1?o D���z��'�X^�	�z�(�&EG�7g���<�HN�2�<�����2������yF2l��Դu(A�9���W��^N��w����&03�ȳ�*�P
��"a�윢VN�9���FeF�Iv�6�rf�"�u	S�t���AC�~�}���u�ı���}�K�B���w����.�ɝ_\�Ty/<���L� ��P g$�~�.7Q��@u&�89�����v\+��Iv9�ɑ ���(+q6[Ċ�wF���'����`Y\�ϝ9�l?�y�n�¼X�3��(͊�}�4���艳��r<&�^I������S�pG΅V+�ieB���=65����\	9y�|˥I���!Z�.�ۃ����%��o�Yİ��kX�ly
y�z��}����E�d�yw�lqQt���{Z7T��f�{K�k��V��=��fmK��a��3
�
�\�Y4-�)���l^�~�+�q�k��C>���mkT�pܚ\����e�aӻ��Mc� �Ȝ>_�ng2�,�cjy�ϜB�%Q�O<���ţ�Ĭ(�B�fW����3���Z�Ex���Sm`����g�����Q���w�Iy���(n�ɩ
v>�&>��������d%r��T:��"��V�"������j���J	�Ḵy��Ҁ4q6�H�$\�^�u_��Pk"�6�Q��F����?�~�ʫ�J�,?�E,����oc��\�^B]L���M�����{o���q}��������8S��R��o�?|�G�E(����񼸶w�6pU��ӓ�x��7��?A��ǴX4���C�_%hʘ�N2.��r��&�+���(7n�QH���Ѭ�5s�|��_x@�o��6>|�=QXմ��D!���5�B�ws��脉߬�r!C3�7%�R�C�|xYb;��r���ʩOl����ǁ��s���?�0�Ϥ&��3!�ӄV�Y>��erƪ�r}��=73�����<�tNM΋G1#!Lq�wQ��.Nc��)l2�Xm����K���i#Ӑx{;����[��Q�%�ŕރ�k�,j�5	f�bq9�DY��.aN6��I���C\�|�7
�&m �O9LN�����������K��8eL�Û\AU���E�s��g��ӗ����;�U�;���?����\W��W��V?����o���������K��}���k[��������|�VSS�|0���������0�"�_�_����З��m�E�Q	\��̕� ��"]"ߨ�(=��"R'��ŹSKx��'P�%��u!����[Z,�M���sx������O��w�����º�Z)`���Q�u-͌ث�R3b3�ؽ,ِ|�l�Ր�%��D�|F�O���H��_���xx�m#���ur4u6J)M8i9)�fN�ܹS8A�w�r�����8%�@�X�����=�X�m�AK��í}\�}Z��0�
��1-1^QNe#M�� �q��5�~���.��"<��mTXw�Z�Y�U�j�*Z*�=V:G�8�əe,�,`o{+�=x�,ve�ܠ֡T&,�u�~-q��/�-qd�Z��~���}��jzL�Ģ���C���»��fG�^�$	g���K�|��b	���4v����';�����7D�u-�2]��ΕJ�+H������>�Uu�$�X��bibVN���	�=����|hV�e]��Y[���&޿tI�R�tU?ev�
�>�q��u�F�s����ѕ�ճԸ5ת�q@��>���c=��y7��oCҤc�Ǆ%94��iH���.bGz��}Rܹ	�2.b$9�s�F�qt���nA*\|���J5��	7�~�($��O��_.�t;k}CQȬN�)�k4�8�@>xb���N㙧G����uԇ=�w���{/��GZ�6�����*�7�B{���� EZ3*� q �0�j)�~Ч�]�����l�P�����eKXh�y ��B�>���MN`zn����vO�軵���e����E��3=� �Bo�d�Z[�p��C�0@%�G��Lqj�~�D��ٚ9r)��Kkj7�q�OI�QR���$>! ���K�(�<�x0+� ݈Xb���p�4C�� 0��0��
���=��k�Q�����1!�6!73-���-��S���#�\@n��MO1
��%�RΕ� ņ��W��{��}}���	���N_6HY������p���g=R�w���}�(��Q���]�Z:7����p�\���e�Ѥ	w��{��]l�2_X���rN���]�ְ��t��@�a��=��e��X��~�a�!�H{�-i��
��SSR�>ĭ���Cf�Fs�z�.��.��	��u��QS���!���jf]]��5�@'�t�4�����h�P�9���E��ryv��?���71/���e|�/�3�dq�L9��I���O�C1�Ô���`A�4�g�t1}jˬyf*j��0����|�q�_��i<����{o�G#�R�ڝ��#�ݨs��NBJ�6�
�5g�aQ����x �<*K&�(K��_�:ב�^�՗���*%�a���(]B��du���3��e�G��w6K�7�L��yi��9��	�zƎ)�J}�w�9�����g����6Ȳ�P4omY&��Y]��-i���9�.�b��	L�O����0\��vq���Ul�%�u��d/s��E	��|�3De���V�c�1j�7�HF��N�fb�r�й[����#�V��
!k�oc���l!�Lf�ZmE�2:3���2l��K�K$�;�jM�͍�V8y�8���3x��왚� va�����0�˄"��(	S��!_H5����<�Iʜ`�3V�p�y�at��=����
������c��0���⎈��U%nUgF��;U��B:׀��~$���r��l�b�7q!;e4��piژ֊�t�6<AR���/m��kL��	�_��}�#ː����P���	C���cg�W���2?��c���vww�/9��wuZ0]R hҊ��m����q���fN,c;������QҤ�z���)E��s1G�KI�&B/��j8`��H���nY��Db��n7�E<�x��54�^Gu�],�y�@��*4���R�IS��>:�U���r��������Bf��u�����s�y��X�2>��;x�wźT0~!T�E8�O���KzB�vF�m;�;ۊt���5�8vs�B���.%ux�/��K6s1_Иs�Q�����v�(\�ո|�*�����N��\7����(�(0$Dl��603Q�C� �U�]Aޛ|ى	���|>��X<6mrSD�bXʶ�ʊ[�)�E[7�@]�t�Z�����q���:��/�!�֟ пe3hFam����y�� �6|�RH��N�K"�kƔ�s�� �䴤�P!�i��.�B	�=����J'�
�s�������<��{�9������/_�����͗0rb����{Or�%��&�2x"Wފ$�q|{O�й�P*hI^B��L&6����.���mӢ��������/ڸo��h�f��4���/����f�nc�M�u]>�j��Y��[���1��8���\��.�#%�ilas�J��v��ƺUl5�&{����䕗p卷1�T�X�>������k�uwwvtV�
�=q��j{n0ron��h����A��R5;=#BzW�W�[���cAZ��f֙�YфM4zd#�#I���p��|A��_xAYϘe톱���?�#
�Е`��|`d�]̣-9�I���:r=�������{�gǍ�x��k��u??��_�޽qNϜ�P�Ag��&N�L��>�szn�&���B�,t	?i7#k2k3
\gK�$Ɂd�^�ãrpɼ	�4�q����Ľ��u/x*t����H� f���� J�,Q�e]˖W����ϳ�>���~X���m�֕dK2EJ�,�3(�D&��Ρj������@��->M`0��Uo�'���aS ���rI�X�i@}K�\��?�ť%i(�r�(\�+�RZ�i�kXRC����
by�i�=<g�\a��Vר��.�ꖸ���E?p�!ꄑbu��M�1٬�۾�t����r*���zc�A{�p/���u���sT�M3u�nʎ�'/���rk�ګ��1�!9e��2tjf�>\,Sj`�Y�.���Z�)k�=i�!'C��Z��1(xy�s��{=T�p%Ɣq+���Yi#B�6FisC&����ͱ&V�.�ϬA������D��!���-���luv|8������rv���dHi:�$l��>�:�yE[At���-��h�|:�N	7z�-%�e*�4)��3���}�����.��F�,���i᭚q'Xt��Rl���|uᱫ�*R��tC�cWu{�h����2�����\�5�[�C^{�D�Ж	XA	MJ4����q㣣b	m'�H\���7��cG��g~%��J��Hk�����������I�F�L���z�N�M���-^��0c��E$�+�v�w^E�"�g��*��%���^��X��|Ꝝ�����k��t��.��7HC���Ҕi�˹��l��a�>�_�W.�R�0B�\�߿(M��|�h����E�������D�w�������a(��08?<l������͎N��6ֳʮ�o!�=�A�FllRh���A����L���a���~��Ɔ�o�F/������ #UX��ε��&cؖ�d�#���"$�i�]fͺ)S:�p�x'�q���ǅ�:���4�y}42:M�wZ>��@��%�����Y�dڴĝo)54^�f]���AwARyA����#a�ģ���e��ƥ`~���a놟qn�]d�A³ �X����� ��ʅ�y��/�����eV+�u�R�*_��Pf�e�dL�&d� |��Y	AN�"g ���K앬P�"Vx�����S���&�#`�8-AQ��]i����Nqnڜc�/�o���A��졃�>ʻ��X�M�J��~ʨ+����뗖��/м�G6ݛ�����r��Jӑ�txt/��/�0{���k}5i_oUi�ӡR���C�vC�3�B��5�m�B�#,pZ�P��	����=0����p}M����cE^�^��=���wj�n����4�^�B�%V�5|����������զ]�i��qg��m�]����T]?�� �j|f޺.:��5P�n'0y~��Đ���|@^�٨ �����:[���+t����v7�c�G	�΂}\�6ph�\�?H޸�Պ�;Y�2�������0���5��e� ��iyp��FXX��>K��ɷ�?�	�sꔜ��!	�PJZ-C��5��.L��znk�c��|��L�P�C��jCh�p`τ��S���(�CQ��ާ��X`���ӣ��b>���AxbM�������M�����{�}�txb�
})�O��SC<ME���s��;g静-�(�����b�ٺ���#�>m��y�������hO��,|�,J���m���u��P��KZq�}qX���	��p;pw��#��Ǡ�������W�abl8�@�#�@A�. ��wߥ�����(��Q�Qa��$��Bj��:]:���q��» �_[���
R4O|����V�6[ j( O��
���`�>=�AG��*+�ӧ?���FFƤ�.(N�x
�ofvV�����M�մu[@��ye��~�����4#���r��@ �nl(P�4�kJ_j�t%A�MWO�]�N�I�=�+Q۸'��r����d����`zQK%^�R�>~�cړ��T/�ެ�|+�!��`$d���i u��>���ɦ�՜�]\\����S���MG���^���Y��k��4�<?�"/�4�O��@��ue^���/��2:T�yjz�|�<��ٝ�V�ϥ��
�}iv��\�ŋ���~[��x������j����Q���E�v��~������FBǈ�Z���j����!%-�,���	�2*7�4�������MS3劥����k�z�[���~rX�7J��FwJ	)��.�~mֈ��e�$V��J��n�>p��A!��������x�T�+�8Q�Ag��S�6WbCao�F\�lŲ���j n�+c�g�kM�*�N([�H§��`bX�r\KӼ�F�G���r���-��jDC��2�aà@.����L����eؒP���K��U8z��P-�y|db{2�Gw���O�A����� ��e��Cf��A��|�~��ӻ�NS��ATK���f=}'qѰP=~���)�4k�*�i�O�^�"X>��p�![�*A��z �̳{��7\���k�Uٜ0퀋 �I/� ߰I���{��	6-'�֠��І��&U
B}�mUp5�%�
��8Jm�m��6��p^������CcaS��k&�y���X���8>k֤V%1a`��M�ؚ�#q��`M�^��lM��32@�5ZY]�k�t=��ˊ�X 9�����1:�	 ��g��a��&F��#�>>>!���o6Ep�i��X=�ȶ[��@�0��$[k��-���I�$� ��C ��M��cwq�*J���34��o��"�e��"�J!�b�9����+�5J��*������T�VOJ\L�L&b���J�K��K��7��4:E �O+#��KB�Fsz��?��:Z���>8��0>�G�u���%Pd0\��00�K�
T��Hq�5�jIɆ��7VjSj+A�k*���b�7+u������֟ӍK�:�6������?a��ۏ���ϱVqsC6�����p�:"�,�ZpQ�d�%��?����{�"�p��F���jÃC��Dl	hv�n�-a�l���zܳ����ߡ�'����#��3O��"�E?�t3r�B
"������e�����=["��ၲ��
�-���S�U��jԈ&|�Dn��¯щq�	LF(&Q(q����n0�*ɦ��w��s 5��lH�{� �)���T�6����m�.b+[Ǵ�	a�Y���n��f`}SgT�QQ���⹣ng�Z�,8��z<uS%ϱ.%Ǿ���Fi}cM�p�n����K�5�b ���{9�+d��ҬS�����g�Br�IY���OӾ��:�&�?wN��[���;��7�̯��m�&���4*L	�1W�fd�(b�<��H���@<i�j�E�\�uMT�E�������y�x�F�ycX����K�J�f�� D�¦C�PQ��Q<q�x3ml�M�������z��g�P����E	=�ý�49<JY �p��{�m�|d���q*���b��4Zdk�C�I�%�fo�@'��,�s��$u�I%���j���o��8�.��ʊ<0���{[8����V�^au�NQrBn�����F0	G�2ipK����z����u"�����K��T����z��c/"��HV ϥ���-�<)��S�?L{z������?���#HԄCR_e�g�Z����4T��s������8az�C�`P;ɬX78�PB��x����˯q���x��{��B0�y��]�R�V�����	%�������B���>:t蠸(h=J21��a*#9����ǁ�������O4��D�V]��u�(��--��X�,��N��#�e�k<����b��J#���
��8��r䵃 Wc6>���:�+:�m�tq���a�椾���k���D2'R^f��¢G#G6N�N�0_Y>��0����$�O�qZ�L y�����~�0��0�'��H1�_>� d2[$u޹�y��p���7�zS��Є!�����n�㷞��I�zU�!j�f�k���zE���kL:�:��I�l�N����,X{q��^J�]�G�n,\Ns�v��U&cV��6����#%p�!��`��G�
	{ �@q�+,&,>�nG��`��i��ŉc]}�l!��NM{�z)�.��y ��偟�1.��}G��P��6�{g���җ�4G{�̍b�P \�yD�.8�d�K!&�d���L� ��dvB,�X@X�$s�kx4�Ry�v��Q,��Xt�k�0��(l\C+��6e�Bc�д����uQ;�C�k<�P�`=;���F��,� J����@��{c/��?� {n�����	~V
a��e65v�_9��Ԓ���\��n'I�7��I�$ۮwF���C{�jF- �����Ϡ�Û���454J+ˋt��E����gqq��Wj,d�����
!\��I���]][�,��pW!�؜ ����@U�JleeU��!���	V�R7l4bk�*/p�O���N҅������KȈ
[�*�D6%�+'E�.�WmN/R�z�����UKf�G�IY��=�Ω������ҿ���a��Z��6��mnm�4
�`l�v� 0��:���3��@蛷{�Q��ٵ4H[]6�����iG���|UEB "e:����q)嵨�v���
wR�"��X���׵tб���
i B���:��<��ZfolC�k�c����Y�����}�{hbx\pc ��v�C�5:}�,=��/yo^oL���i[�т&Ev�l�kN�W�x�M�w�#���i��}�a�?��wi�7���������{A��1�x�/��� ��9w�9](�XA�fS���
����aS�CDTM���������E_�E����Z�C��ꛏ=F������%z�����~O
~�M7�$�
}���7:�.jS � E_Y+�i�_��*mlJ� ZXvL�u풮���q��g"�v=��GQ�r��C�xPx�v)�hX2���|!/�F�1�H�]����W�X\*���J�i�Dh���G�'�g�v��/�Ɔѿۺ! �z2=2Z��B�|*+ô0�U~v/����/�8�ɱi���E�)}�V�R�)���g�)�~��ac�X�r��_�!}�����r
w�hA �Nm���>�'�\��AS����u��/������k&�7�MeMmZ�X,I�)rb�I!0�;��S��ہ��A^�~A�hV����9�T�@<r�� ���ӗ��ie�J�^����vCWVf���汅�{$��Q�ي�]�1!��-�2EBH��1�N�[�U՘�:&9�D���Vι��I鷜�3)��_x��_8��ܔ���»�� /S'hN�ǂg�3KعS��b�Jʴ�����'/�^!�vD��'��8ͯ%��i~~=`���P���e�B�r��eY�����W%�ڛo�%6�>A�X��C��L�}�,��@PIk&�w�|��6o��{��?<K��-s���(M��d � � 
��Ȑt�í�uC�h}�˗���!��#�{8*� <p/q��J�1?W�5Ů\��-r4t���G?��JI�
���G-_a���0`����X^�3���,�[kR��`o�~�|>-9 �eDP�v��V+[��D�Q�CI���xl�g��c���a�7wN+��Jn��r�y�C��KT�(
�P�<$�ӼX�zT�W2�t{�];�ki�q�lvp����]ή����1EE������idhi�4"x�B��Z���f��}��?@��W��_��=��亿��o�M7�$�|����ǿ�o^����q�"^zUQgE�u��|��ZP��+�ᰪ���11�Cvc�F`�0�Ɵ]g�yj�ʀQ��+�HK\&��t�V�QC� n%�� ��.[�\�b<\H Ƣ��y���f$���	��i�\�.�=�Z�3>�S�]TL�X��laӤ$(��ma���{�$ `B���FH�<��l�*dKc|i���1�(:$(�]W�~�4���Ƙ;�Aq�y*b5��K�
�+���8�˕K^"�)^o4�OKb���$Q����
m��J��e[Tk��eP����L.�=hB2���  >j��� �" ���t�X����t$�� �b���-�!�!nW\c����qi��1��O?��ɪ�����݇����'�l�����zѷ[bE��L�M�c�|��V譏��<�Ŋ-��"~?yA
k�mS���hY�q��T������Y۳�� �B/�s�V���%D~��I 4L1�)�xp�n�WI�#G�ȢA��B�7WTkbM�$�����a�1��ґ���Ȱ��ͬ.�����)�h�bU�� eQ�!(c���f	Z�XU,�$B(JX:��S'L�H�'����YK���B���[Qʲ�9E�~G�e#˘�1�i�pJ�g�2I�>�Hۚ��X5-U�:{U۱�v󾮠�Z��=��J����zDw�����p
�0 ��g��`��؁=Sl!=�ܝwK�����"�}�!�~���ǂp���w��n��f��W����lq$|�;��@m�ͮ��~�0��7��y��@B|׏>����ߑ6�g>�����/=�̳"T����ѽߔL���5D �f�h�1(�õ�T3�=�Hr���f6��C�LlÂ
��U�o�-�7}�N�q���?��=�,��������D��960ܢGv`(j����:^����I&�(�Ǣ��*�}�k\N7Q�ý�g�\j���
x\+K���鬰��R��j�Q�]�f­FS4N��������t������G띅ngrF�"�d���G!h2��{

&r�p�UG�=<�w��^}�U�_�����7�~K���_Ϝ?Cn8 �t� �B�p��;�y�(�㛶��+���0*+HG�o�6�9AR��$��M���������e����b��5�Fg��Ǆ��m���K�}�����$���Ύ�@� =m�j,��-�Ϸ�׮W���}�A�ew/����U]`�)��g�6��E}��e12�gm��@�Y��v��HP�Cj�Zd���{b6�zzAb�;��;�5�_�p��n+0e�)�
� +-|��Y��VY91���q���R9ÿ��>���Z�0��x���i6^/[��N�(+�k�߂���j�ٺ�8G;FF}ɦO}��]Z�gY!�����C���å�?u}���P�KG���"��"@X�[>{��ߐ8�ыt��4� ����y3G�ΛiS�T�ma��K�Xw���$u௠-��?I��"z-��B��`��0wӺXp��>��:ʷmf�8N�BI\7��H�(���O�U���iܵnG��g��?��^ݢ�lJ81�\o�ۏ5�A>����"�,8:a��n؉m��I���H�3�++�Jw&��IKeP��0�Y�����u$�be�7�Z�ap:�M+8�S��:f%^�8���d4k�Eu���=`.�$�"�8p=]�(/�p���v��ϳ-#b)J��b�+�(n-�`�(����hB?ã�Cb%0�7�֕$]����;Ƴ��V�ͷަo����z�����̴����������ij�>��o_��-\!��Fh�YH��v0� �q�,�'"� �&@o��s,�&P�s��hn�wt���'f�b�1��M]��V�	��V��M�KYȱcG%1�&lX���1I�����5C���*�q���le�H���7�'+�Vo4)�M�p8� ��#+�I���ЎQ�v�1q�/�(!����Pb�/�d;��F�;⦰��o7�m{q��xs;�!-BkK�%4�<<��d��գG,��f��(ܛ��];�$o{�k=�,����M��ޯ]_ۤ��ֹ��OC���ԩS����N�f����H��-�سΉ���߼L�gWu��f�L.�v��P�7���v `���������m�[��erT+�ECj�B��$���Б�{��n�}ô<=K�|[�n�j5�m�!'����m�',2z�c�pN8݊��"B��;�U��B9Y1�X>I)����B6��D�[,��*���\��C�������_������%�K�����2�q�G��QM���[���t4�:a�v�Mm�Fy��N����O^H��R��K���I�~���/��� aM���_$p����8�N�=.--��_�l2>e9�x�h�^x� �4;���/Q�ɮ��z�^o5(�E#�*e�M��/D�x^;�UI��P��th��׾N���ߦ�t�;{��>�;z������6�(�����.h׽{�H�)>�R�l��ɑYX|w&�	4�=��N�#�>B�o��-t���������
[�:���	�uJa/��*��W���v�Ƚu�>�A�F6���Z\ϱ[�;y��l[��,D�r��Q 
�(�d�4yعѝa���,s%?����Ҁ9�u�d}U�	;O�XQ��v)70L!yx��wѽ�G{��H<��;����K�/]�x�$^Q�'a1�S��#�/�uǀ�Ʃ�2����'�S�N��)���iJ���'�	��&�uZ�X���:���i�c�j]��l./B�7��,S��Ij8'���`��0Uꂇ�ʹ��鑘�)R)�ۃ���*�'�|�˗/^b���Xm�H�keT|�����@�fͲ��Xw)�)]mQ���|.#�,p151�BlR��W���8n:A�
�y9�l�Q�B��un�� �b�X�
�7�L�h}cU�����&�m�n&����d����ɦ�뱛_�@q����&f@�#U_��T�%�W!x2��c�y��œ�%b��N���M&�d�n�g�#��f�CS�H��d-���6������>p?=��o���o����4W?p��YQ��O~�Sz��'��1o�����-:�5-�}��`b� 0*���c���$6��7.�����-� ������^y�ה��ed+!�����!6Â��yvv���h��-�S.��C�B�,-\Nhq���#2���h$�b�tH���~ ��!�U���uL���#�p5R���j~@�+��95Ņ�q������z�/i�]"7�0ۄש��v(] he�d�4��z)3�z��8�J��U�M�*۲	��a9R�H�	_P�Z
H�pw:Wн�nj��&>�m����	7[�}��GY{Wj���O�Gt���iy}���E>�k>99I}=�����T���/A��5~e�0X�1��'�]�3q�k&���l'�f�I���@�[aˁM�8HnH^�S�X�����
?�|=�BCMɼA�
m���*��ti8�\~Fl���dJ�FS����,-,,����ژ��1���q,[�h���~}o�}����ޢ��e�S=v��u�X�ޖG�fi��KH�Z�ڭ�|W)�����p(��Y;��x�����z;�� ���.`�_kk5�N6k������ш����m��3�{;�e`��1P�1��?h���p6/�qv�hALcW�ƺ��X�7�K�D��'�$W"�V�ڽ���������t`�q1��'�J��nd�GX�?�����/���x��W(����1΁2�V��:c>���[Bё��ծ���
����� �hTmHp�7<L�=v+9�5:����Ί�AX��ig�죱���61��J���xyI�%-7h��պ$פB�!ö* �) 'w�fM������g���i��B�u.���Ћl�k�eID�&3>J�c�D�[T[.�$�m���vty��9 Ed�/�9���@�����Y�ik$�pf���0�����\����bE-���"�R쨋	���n�k�P5�N
60��д��
��J�u]�e�H�������D�������g<J9����|�N�9�Tn�B�o����#G��.�!���N�)�i{[���L�/�Jye��W��-ބ�*�'�',Fh�4Q����l�s�m���=��ݟ���9����O~�;I(�8����F�n�3Ǿ�\�ag�p޶�6Dkۍa����c?BS��f�F?}�i���P�X�z+�����c46>A!k��VM2�.��~��c����ژl=
��2`��`���5�wm���5P�]Sn"Sm�����Wz&A#VoD�����M�T���q����3q�vح�f4$��$Wo�|�Ԍ�Ki��W�g�)����e�%2���?RPQw�����Xf�t�LXugW;'o�(�?�B���h⍵EI.rH��O���& �V��z;��x��sō������Xɳ��ͷ�� }�dm�:��V��N
�83+���k,��	D���H�2���
E�j��E<Js��P�>�xd��A�r,�K�[����in}����]3W
��`13l|�z�|��ϋ��ä��{��1l�6���[v���'SV�䛭V��_u��PxZόqC��*�^��,h2"Ԉ����g({� `�V{��;Ӹƍ�MCι�	���*� �9�?�yG <�S]%���t�`/B��i�Ӥx�P��n�u��N��/�
E��E�b��v��t��-�Μ�� �PEY��v]L-�e�5�������OPǀ�]���V�o��nqm����3T�`M��Z�]�6h�Y �f9fi����,���AĞP��6�}��t��Q��R�q������n�L\(ϋ�\NQh=sõ��w�}�9Ф�FN�7Cr"��2�LN'���[�Z�J�z�����(��
ҢvU�- ��T�/Iɤ��WD���95���T�Q��[~<^d�e��I�&$�B�v�����Lѽ���޸�	%ߗ�2$P�n�/,�PFp�1�ٍ���1�}��-cu AG���ͷB��� �uqࡣ[&���656KT�[�啕(��\T�w;�J��*%5E}�F����L�W�J��;�ދ���m�����2�h�P�7e��h�n�x��aK^iK
�!m�)�Eɠ���՟�0)���vZSmv�&+C@q��t}�v%(	-�}�_����E�Y�GGtt<������i��`��=M�cp��E�X�8C�C)��I����L�G{ȍ�)�T ]��*DG߃k��?~��u��J>�RB��94����tV���R�PJt]8W����~���ZzWMW�"��G�*���͑^����bڜ�Ȁ��O�օ96�u�,�|�}�5#�&p_$y�2%S��d� V�9P��S��Y��� �k������KK��1*z3 O�7���p,�_/`+�r��YN��i_�0Ф)L��C��/��PG��l)vm�څ�M�&���,]G��6;q�kb@<d׸X�I��D"3�k���_�Jɬ��z9i�Ɵg��1׶ͮEh�tJ]�\5?�׸��/ެj_bP�B���G�8Q���Et;^�Ͱ��.V�XD��o\]$۴DE��$�õZ� �=���ިѻ�# ��}�R���N
R#��܅s������Fm���Zǹ�lgD i&��C�E�=�ų��&�Yk�������b�q���:�ZE�a_��hX�(�p~�U�q��c�)��5�G� �N�`�\!O��
*
���Z�Y��hV���^de���EƦA#5мj^�*�U��CQ�7�f!\j�yi>���'�H�s!��<q��(E��%��v�����ҝ}�֑l����&��H�m�i��� �I����sM̔L�d�cG��m����L��m�N� ���0�8G2K������Ա������D�ۆa��&���Dy��x&>$Z^}�u��/~���/� �ʦ#�@0`�3�~�8����>�4����S����b������R��n��J	�o�RȮf.%���������O��0�l���ӧ����J�PPk=׿��)����鏿� �[>���#��o^��� [��W7������~M�?�(��O�{�w����2=��CR��;�K_{�U��׿N�Ѧs�/г����5�� a�lLY���Zˊ<�0�u�׉�n�|um�DG�]K+4�o:%�����l/�t���d�������:�d��z�
��Ɉd$�܊-����kv��DK_�\`���?z��[}:M�ؑ��m/S�z6�9�V�FE��+�?��@z�Ql���D���on_�F|�5�n�����a�.��y>!uDA��K��]9�^�Q�������uZ�m�H�(����F\��(����߽��٪���
�z�8�P���9m!7�8�W�Z�g��g��Yz���\���Z	k��
i�-�(���O�N3�u*eE�FG
�D_^����DB�Z��j�${&���ҍѫ��}��]\*k��8�O T�A�f�<s�K���4�TW;�����{f��l*^����v�I�/�����u��8���C�H�5����1(1�t��kM��o����yz������3Z㵺���|�z��7���^W(y�+�C�$,lG�%����>8��HG�U�X�kf͎��t��ꕃ��7�ϖ�+��7_�7?~W\�jY���K3���P:O/����g���}�n��;�Kgf�}��zGF(���N��o�"�G�}���ӹ�%:5}�n������WC���~�?觿��J�8=MMve���?~h)�����d�d�O�IM�4��.�����{Me�q�w�Mlw��QC��!����q�ZRQ7��kJ�HF�D�L�hf�&�:%kp�ﮫr�z:������V��9�~�t�G�Ld�0��1ֳk�[kD��b���i�mK��1�uk��5���EF�ˏ��p��1}��>0Lt�m�����_�ͷ�LKs�t���(l��8t`x��x���?� ���?ѳ/<O�ˋ�9	6(٩����R��k��|t{�����}T��S��TqYC��J�X)ʆI�î���+��tu���6��rqc���_�����H�N��%��e�@�*�n���@�Y��s4��?��Hu��gJEz���h�����Lk��Z�l�0��69h�{F��c7�D�X���`���֘ ��v݄&5-x���X�g��+��*u��������S�����ь�M�_2���@�쨌�J{��G5J[���/�Y�IڔJ��G��T��L}Ԃ���΄��Gl��O�1�C��k� �}B?>�C�'/1��y�}�r��t��#t��Ӈ� ܆PLX��o���q���H���y:��{tiq���ҳ����m�|[�ON4\mt�{���xl?�d�`�}sV�ʹ�e�C�Q�q(����Ix�t���:����|_/ͱ@����V�*�d�tae�J+E����m�E�f��
��]S�tu���
Ο�$����Q`]�2���# ~ 	��ײ���(��>���B��`ɱ�hSV��d��Po^��8}E�ȧ;!��F�zޡ��wgK��ɰ���C��e����"��iu�McF7�}ϋ�W��ݻ�4�·�h�,�@��~������ Y��~���8:�e�2��Jr�]��Z`0�����+]��&7������i�OPap�n�� �g���Qﺂ���4��Z.�����;��u��g	�\M���P'�S�RWMӛwo�Z�-I��$u�34:����Q��x�TU�O:���|#�w�0T�nP	�����e�!�A��������+sRS򑍅g��kQ��0�E̳�Q-n���� ����{4�.aB�#B'` �5��&L�#��-nZܦ�Mb�����VXKt���{�Xi-���1�+�'��N��C��'��(�[�)��o�Z:�Y�'�+(b��O���a�M����]��w���b�w�ʚ�2��T
�����8�HG��nx`���[\tu�� y(�o�2��n�L�k�t�m�H�/�v��N$�{W�y1J���,Ej�&�I��qP
 � ������	�
���:h�Ҩ���ݓ�=��IKΕ����~A�������i�o����1�F�L��*�lU�$�����U�	>���*j}^��-����1�o}e�z��OК�BC��.-/HWJ`���Տ�/C+����9��K=�'�����.|G�*�˫T�_�%�ǁt���f�(����ٞ�P�3����Lc6	��IX=k]�rVeZ��AX�9�q�`������{X�<��+������Jg�b�!�G��
��@��ִ�R�XIey�+�
�5�|)�:GY$R�B=LĠ/��"Qnm��S����a�T	L�9�&h;y0���-V�N���m=�*��8�۬��]�V\+��4��A��uϲQ��J{��b9-�,4i۸������z��a��S���u4���� �
�(���p������"�0m�[��P�>�1���p7K����ej�6���{xa
fr���=�בV�H&��p�H� a�>Ī�۔�n:J%�^3��V��8Z��MZ�[��ł���G�V�s̚V�#��2�\-V)������Hz�u"N��Y�q��	w�Ԙ�s�ڕ��E�C٘:'(�_�Z���� :9�ý[:.u[=�dE�g!���.%IN��&��Zd�s�kAa:e�&��q�Vd]5
Ot�l��C�A,�E�(�Ï~���>Q4��M�%���<��#��]_��/���j��R��L��3��q��FY�$�c���f(�2��ղL����DKz!���HC���ˋˬMS�30HMv/�a�є�I6��PX\7�ץ�'`umc]�y�*�������D.�t����.2M�Mw�GQ�d�Ӽ�f���+#O���}��u��t�4w�5w�ߗ�x���]^�סP� iA1�h��8���L� Oqm[���ٸ�nd�ق8'm���;�r��p�i�Q�A�Z��Y�H�bE��8��O�T���;q�:-�$t ��@o:˛��qo�ֺ��_��T�)�v�[m�5���Mx)���@�~S��p-(��+VA�Q��'ߢ�ﺃ����K|Q,�.�enT�@tx�����,��d���f&ɖvw��w��j����c�P��$1�r��:W�GI�T�l*�z��¥��P�RȂ6
CepI	��q��K�E

}��i�pǦ�]<:9Ac{�TpUX�[%0-HϮu���F�K�3�JX  �)p�.���	ZF������(��?��*	�
�Ƌ��k��3&ntik�B�[|�د�A�(k�S�b̡����7�%��6�ǝ+���pB%�V�.���M�LQ#D�4'���a�	�:g�+�NʻN���L�����ޛ����S ײ|ɘo7o�ۛ�L�k�S��X���:[�N�pezq�����"�_��I��3<��I-��O��~���r�pgk��6۟�j̺���$K� �a�d��.L���3^J�M�5\�|�̶����� ��^���.��.��I��u�fe����<���"��ϟb�N��1����JG���0-q|�AQ��q�}��/Z�Ҭ ���M�Z��t--����1��!����lJ�L��-�),x��06�0��?6ѣ�crˋ3�0=�B�����a'M͙����&����M��Ic�[A�%��1F
����D�l���d<�؅źB(�tx�Zh��	-�Q3� �K�}��P�afmk�^���xCC�%`Z���1����|�{  $ s�Ҩ�k&ѣ| ����7���	kl)ü2y�����(U����8�-��@�9�/�ϕy/�� b��g�{�S4��D�~�U��؍4<8�nyZp�~��Й3gu�π1.r��%�K�:lfNږH�O?�gaI�����=�<6:RZ桺�X�m��$M˳Ygs�C&qdD�/dB���M"�?��qZf�gA����I�����5ZY_�02��1�
C�4��Lё}�)ñۅ��قV�JU�:L�F�0Ἰ�xl,v���a[�j(�2
X�Y�J~����aA�ѥ���ij�6pM>L��_Z)R�TVViXꌛ��x��x;����")A����\�j�f��Ѭ���G���MZ߳G����k�v��BɆ�9
l9Cʡ�x��#�
b�x/⢙b�$%m�52��4�1�vԸn��:�;w&	�e�Z�g����1#��vQ��{`�}��W�[	� <��\%ل�C�����6�.|]�5�np������2��d�}�/l"Л�C�����fT�F�"�!V��A�(0/�B~Հ�ע�t�`�d$�֗륑��g�X7�CS+�f��Ǜ��#_x��r�g��;�G?�� �"C���NMv�Q��36A�l�S��c�#�fer�����Hl�i�^a�J\��Q�F��=?+
��Avis����l�|���G�$��y|��g��V{R�9C�h?��*��.����K8���#��趱9����G���J	e[.*�'@����� i���Q�L�Bv�Z�0n�K�������ez#!�P�-�Rv�.v�Ң���Rº�}�3�vk���SkE��e�N�U2X�{SǗ��g�f�A{&&顇�F7="���o������ V�I`Y.���N��!�B���"���]�����a~�2l��@T�50-C�C�T�O�o�͟mI��Dh��6�2:�[ӆK�T�"�ی�t�z��������9*Wˢ�2��{xC�a��� ��]�n�Ϝ��z-*4�����7�ًg�ݳR��ibj�n��VJ��-бc7ѝw�M�9M?��S����d�6"# 6%�l�����/fyqV��(�gS=�wb?e٢�M_�"p�7:��9�r�|�wF��T\� ؙ�QjJ�fM�&�^$L�e�xp�`� �(�3� ��28j>hN�-��� =%�?aH�)x�2��F8C�90���mUv��2�6.R	HZ6[+6�b�Rt�gt� J�"X$�"�'�f�  멥]�W�L�X`���
���JHD��C	��=������<}��������Żo��z�z��稱� �G����\�U-��ƶ��$��1�0���P)���I�&>���4K`.��Z]U�\�]7-=8��6Mv�I˚bS�p?�qL5A�l�`g ���7�὇�U��/��gG�t��*�sTߪH\x`�>^�:>�O�d�p���_���N��x�ei���N�� [4��LS��_�p��ert�VWh�]a,(�4�Y���S�����s�X٢��7��֣�Z���e[$p)0�����+7��f2�1����5�2
������B +�$	x�n��T�
�~��e�!���yD3�/��p�\
V�  ����3
�x�B��x�Z��i <G�kbф����.��#�� 7�7��Y���q�H�,I�I(�!��[�@�L�3��@�H�Aʪ�j�BF�����{fqNB�4!�0����O�w?���?�2+ԁ�^:�G��v�z3t~钬���=p�����+�T�brGj����-_8Sd��ڹ�Z�-��^�懄a��RU\�P(�5���#y~7���������Jm7��|�����+�-�~0���f���`��%j�CMcsd���� y\О�����C�uH�.���X��@�%���a�YF{'z���_:�Y��}h|p��g��R>W��(k�^��._�LK��  ����Zj�u��	�
B�qM�h+6։�=g�e�]3o��6y�2"�"����U�R����Ѣg�~�@�����Kh� hGB�m�m̷��uď��ynda��� ���Iͭ�M��؇5���0��h��?{b�B]#Q�$W�R���7����AM>���	z�S��G�I�Cct����ď�������J��r�����`� 
}ŕu�׆����t��RQ�^0�ln�Es�����%I�;��h�.&6��"�o۟C2���G��O5׊���5�l(���Z�؝��(��Ac#(60�=`�k@��	��]�f�J��:U�l=�M�qO(�{l�2,�%4"��e�Y�ĺ��4�Ó���P^^��f����pgX���Kl��\�V�Z9�h8%�t��<���ḿ�J��x�k�Q2�!�b�QJ���;P��*E�� �2��T�PĘ��R��'!lZ^qdV�Ё%�����d>@��a��N�8>i�B�y�zTC�cJ���*QXFĀs�G���9~n�b�ڡݲ�+q̷Y*�ĺ���1k��	�`������|�˞C�u�%^Y[�W4�R����ߧ��o� .���}��м�����9,�E��n�e��\	]��^fiӹ"��-0�4�����[��Ʀ���H8��(aA���E5]S��e��R����WbauY����=F�=y�x�����K\��bUx�Ml}q�.�>MٌG�yZ`�������:33Me���{�00(�/�� J���������Ÿ:�@k�KT�@�,$�M��>��2M�c!���@�\M �a���P4��K�yjM�ckG	�P\<6�s~aA\J��	b���##B��+�'�du2@��Aȶ���zT_Ҭ�/Y:/	F�Δ$��P>LYĘX��f=�(V'u3���$�v�l]�X	�kP�r�=D�nfs5�Y���yۄ���^ľ���H�.hO�K���*���`ҥ��;*-f�|}�{hq}���^�b�'5�)q����w$��NGs�W>��.�<V�ڴ�b��=,�M�@f0!j�@R�m�8@2O-�RG����5)Y@h
�D�j�����%���7-2��mӳ3�Q�w"1#��-��o��U���#���ُ��W���r�y�tB"���Ğ=t���tǧ�/�K��-�ɾz���$�K�i��r��+�ԄAc?>��iǈ�T�f��I�z��Ao��f�����V9̒��2aъǬD6��L(hs�����cj�����Cr�����`��2k�l]�g/+�y�%�����K��@#���0U���l� J�K� ��D;��$�7�ձ�(�;Y*�E�Ԉ��/�E���fe4+�͡7�-�W�צt'�;��c�Ѥ��L�O	�^�[_g�� ���r��+��]���f�D�M���1z���hdh��9A�><%��@H���Ȯ��LR�&�t�,�t��I�vj���~$��0:��w�c�8ts�n�예f̄ٔY??�l�ҎJct�)��`�W����Qތ�/���\ ��@��-que���Ja�N��t��.���X����R7�|s�m�����Ka�����9llUh��yp��ö,��zV��KTj�b�kb]�`[q܃4.���(�lS�v=�5�$^B;���I�;��փ�"�{�d[	��$�+X-�L-�[������0	���0R�|ϔ���ݡ9�r�L���ʛn��#�#tϧ?#��^���D��&ܻmQq�+�VD�uiS��ޛ���K��I�+�^� u�������?��rN���Mz��W����t��ҟ�ٷi|����SbJ�v�l�;�u�X;�����DQ�c�H�A�$��)�ˎ����]�7�`t�nh)/�9��v�����ej9f��xB��XVL?��-e�O15��Luh\�IUϡ��t��;�Ḋ�� ���}!����5��l�"[���4eY���Ws��OS�o{G&٥.Koi��e�/�����_��YT"��5�{`qN$3�j������?4^�o��
�p�P�{�\�fUBДd��'&�{��i՝�@����.z�X���'��A�҆�W(����SPu#X�h��K�"�W���*��Am�����@>G�n8D�l�C3�4Ѹ\�)uM��|��׉�ˁ8����U��+k���%z�(+�'J�����J���g.�+�ߋ/��5G�}�B���ϟ����U��GƤ��ѓO=-����#��J"�.�?]n����(�e���Zy��6-g���QE�wu=��84���w�AGo<,��/���"�0���!�8*��p���bŐ�aF_�6��*M��$�҅[�,57ۂ�����rYP�zz{�"���Wت�q̆5�q^Lٮ�/j���&?�1b>���)�,�Yap�H��͵\��1)~W��\o�c@":�6�*%
���-�ݜ^g�B��B�W8A3�V�3�+B$I������/ h��K�0��e&IH�cݞ�잼��4��|᪰y��,y��Q6q'\�٬dבM\][�UV&�ϝeu�P�u���4{�΋���Ӟ���N=Ŋ��=�Ir=���e.��h-ca-޵|�f������S�C'�$ɭ���~��kR֑�I(\Sӵ8�v��� %��<� 0��o2��a��H�붆�ɐEC' �I��$�.�{�Ņ/�(���#�?@�}�!��]�Y�O����['���<�%����w�I'�Kg�R?މc7���2�t�5��<G����L;t�?Ӟ��"��*���۬�ot��^�����K2������H��><8,�3s��VW�Y�t�$��w���^���M8p��!L�`-Иm������r���C4��ҥZ+�E �:�â�)�_S �������ѱa����2E�#mP�r�A���o���ƺ֚B#(;1�}�_N��1Uq1��8T�9��]t>!�����
0�q��7L/����W�vk����i,�*T����*vA!�c#���/Ub�'��g�d5�_4�^J[��^�N���}�7s�$V{c�]�|O�6 ��LQ��>���b�����xZ����XY[����Q���7���
���q��=�<��-�#qw�|qv2�P'��a��QH�D���35ح��6z>�ѓ�M��w����ҭS{���Aa�H��`�|����:H��CGD�Ne4\�{��4ah���ቧ���gm��F[_� s(��c�5�S�����ڭs@��p��ahÍ↌!����5Z-���M�b�������{��<-1^#��xP[t�Y_�SU �"kvُ����2�9��][+�:`�����c��O�K��(�:Ej��x�<��!m]�mfج�Ag$ �k� IaGvкw�i	�r/����0�%A!S㳼����������v��M˔FB#��	$���~�r�ճψ �d;\���&Y�$���9���,�%ԆS�ԧ˛EI�a|wLߴM�uh�I��g/
��z�k�$cp�):�-�-�)���6��FCa���8�&��2�Q4��
Y#����r�����4D;��}�п�(ў�A�75I˫t��З������/�'d%y�l���.�_��W>~�.�-��R�!���4Hy�WYSi�A�k��a-��JQ�i�V�Ae4I��	1�jF'(�+==�qz��ݔ����-��V�ִX���Y��� �Y���kh�$3�[Qi����k��o��̏@�2�]�������@�ۥ���!I�߂M�I���}���,0����W�(훸1e�=�!ȝG���b�e`a+2��JA�`�����Qܙ�v�
��\� H�#$iv��e+Y�}UaO��)��Z=luY�����p$�W�Q1o��)zf�4�n#qb��%�����/꩹����uTt�H�j�
x_ђ�9	H=}T�GER��۬��o��V�]��jk��Mj9Y8��?G�[ilp�zXHW�luͪ"[�Yf�*-����k �NI�T���Q��qd`�Zl�A���K���:��0���]�8�eرq��x����A����G[? Qژ_�*_7,��������������V;Z_�ذ|���n�����c��Ӕ8Z �I���)��A��}S���5m`��a �lI��40�e���=/��۩[�_�c�3�Z���w�L�Ȝ"+4ԀA�Փ����ܶu�������]/M~6-��='na/ǣ��j�X誎���kn��N;�K���B��c�4��=�ݫC��1�
n�� �J�$Z��|_M����m@������Rm:��ƀj�4nV�"|��ai��Ą�P��P�e�Uh��J..��ři�Zǆ�5��k7U�����(J�,�����4><F+K����)n>��=��k�43=��K�6�f ��G0a�Bb����� �j��ϫ����D�u�v�%�l��#�5F���}���(���Q�!0�����N�B��G`� �B<T)�$*���7(b&�F�Cy	�j�턀hy!I�����S��|d�+^Ӟ\A؊e�5H`Rc�1�:���� u���;�)�:���~2\���Uד���xU�,����>�ϣ�ԑ}�Pe��#��\����@%�Ď;B{�N� �G�_ڤ�Z�V��y��uZ�nR��?o��f)��v[$G�g�*��
�?B�;�.���b���Џ�����:QF?�Z7\�jieSj?>PZ�^%��X��O�g�h��I+����$c�͗��d᫈k��6/����y�=��h�3rm��-M1�xA]jA������a���D�7�4
�h�i���t�,��S�]��oh���Uƽ	�	Z���@Y��W8���wz�3�4�"�n|���sK�(VDc�t;�<Q.��t�[�*w�u-a�J�-)Bò�r�844��݂�B��!��b#�|��2l��|�������T�ޠ��n���&�|�q�1�-K��h��ktt(�rxX�t�%��������4)�XI_k[Q���Y���W$��gtX:�NN�P�i$�����F����>

��;�Ɗ�w-�&�E-p��nxh�C�&��,��(�:�TҒtL���e\.O�} �Z�1��M�:\�L�/�BwN����4]�r��&�3�������c���g��ť˗h��A��S�'M{�OQu �xE�%�7�Q'R!6��5�11>.=��K�R�!�����4k��W.KRd.Ҫ��,��ўG��~�����_���-�8:�lm����XX��ڤ4l]�y��I	����u�����a�y��R)G����2��\x�R1��b�P��k��t��5��8`�Tf4�\�)�،�n��2bTa��	��B�
b�&+�nx*ɽ�ﮣ����j��$�ȓ�}��P�<����9�ZX�S����S� �`�6��0����p?�p�F�YY���e�b�q%�D�y�G�,ҠtăWi�N�t�����4�� ����f>���-VG4W�%�����GQJ�~�r�	r�T�[�{�����S�OYdk�����eZ���/>�w\؏J+�J[�	��ܐf]�p�< ݌�R�χL���!&d��@3���t�Գ�B	��ρZ����U� ��a�8�_�7�A�����ռ9 ��neQ��h���%S���vx�$�l���8��N�!4�~P�ǎS٤���;7|��l���$)�I��$8���V�DM�S=;V�cǙ�&�*���������T���*.--��̌Xyt��D;^#i^;���4�I���n>N_���8��}i��--�ޛ�z�>���d�:�q���@�L����ۏ�C�G����c�F~7 `�>7��tt�B�?4�.b)�t`�l��c��B괐��k�K���t%{��B!���C��dC*��h�e�S ]jq��hi����P-������xo#J� �5�\�2�r�
� �6mCdo̻'��!È���(��7iaiE\M$} A����&i\��ǛDO��Ӕ��k�mQmqU\I���U֤�� ��f�c�w�^�{`�L~l�m���,��f��ΌoI!�����g!��&�z#�<��lH���-sǟׅ�B5�rԷM��N����́�"����a7��&��h��X��`�Դ�f��6�"��ϻ:�b:�hD�fi��T� W9�����P@ #P�45��x��,�=��p�x�w��)���}�������i��|��&�n=q+���{EV�z����_<M�9#q���V�-�ޤ�C��Ʃ�o�řE��Y��h5Vas��)�WזkH_B'4��� *\
�f�_�N�!�	���9�w�lkA_eғ�,��V�&�yO� �P�?�����,�O��^Le��iV���0���{A���7r�E&-�4�n�߷_:h�X��[۴�i[i���N�c��MJWx��DV�(�V��c�;n����[�ӗ������a�b��?��_}�^}�U��U��Ν�e�!�#f�_���ˡ����!t�+C���"�b7F���]�oq�E�n$|�1���5��LbH3��q�[��P�W�:��Y��X���������gP*�D!l��1h�UV2]`�룏>B��Cc��t��9:��iZYZ�M��lE����bbb��?Aw�q������ѕ�Y�nо�96n���	:8>H}�<]����bW�丒��.���7?<ǤF���)>��Nx��H�g_�F�!���+�·�x�i�ý}�x��J�.�='��T:/.)`%Zz薩�W�}�N��^��K���~H�g�蕄��w������gR�Fɣscjl�$/���D↔����±~��E*�&4����i�QR#A%j�lQ/F��}lU�ԟ)��H��c��_}�/i�ԔdӀ�<7?'��|(z#}>:6F?�MZfw��S��
k\��֭�y�ê��0V�A��|bZ�_�
(��;t�ۺ�m�֒���%d(<�v�&׀FjЅD�S�5����B��)<��c�8S,P��ibW�m�X�fq������g&0<[��/���l(������+���ޗ&�+���qI� N�?s�<=}����r~�3��7����gt��Y����}�7ܤ��!f��ë��yZ\-�S��n�&����X�dc��wD
�F����9]Kdc��Ò��/�N@Cܱ��@��=9��?D�y�1�UX���5v�8�6����enb�^d���2}��-4ܟ�����u��M�o[>v��hkޤw�F�ib|���yE�F��η��O��sJ=�JM��T*���%���\���&���´-P�o:z#?������O$��vŃbPv� /���/߇�[\g˻Yb�t�4
���,���۴��"}�m�M�$,^�Z���"�
�J�	`�+1Q#��������Ayɐ?N�[�߻�/�#0�O6��:aK��{����#f���h��bo��
����F�L7	cGJ#���� Lh̲' \ J��ߖ�Z]]�����( ��2
��4�c���2���{�oj}��Wz�]�w��mɴ@d������%�u&x2�/�}WW{����t0�h$��bGڙ	�J�����������M�FnG͌�#�t A� �F�F��6U]�W=�2�|߽7_V��&���W�e�{���w���rx�(	�j�o��b��B5a���V��5Z�Hl��V�5S�x]�p���T��1� .%�
0qH0���.}�'N���|Z��̃�}Y)j�~gN~R"hq�~&%��Ui��8<2���l^��~����3�? ��y"��%��i�*��>d5�����'�_�V�F)��LNHo�]�����$?�g2s��i��@�����E�R7���)	�c'�����//���Ү	� ��m�l�*���`��!�)-aP�����H�q]] Wȼ\�I`N�e�DFH��y+�K5�N�J"Io ���ꖐɄ�R}$��L"W�s�4fM�|˯i��m���T���|��"��}R�ܻT�ℍ�Fv ���k1ڕ_h}�� �02�!��$8k�2(�f<��h(I陁p�K��/Y~S���.��`mj�/?��2�{�յ/R�k�oߺ�gs]׻]������~w@>8��\;C:�R��s�$љ����b^.��UDoch>LD2!v?�ߝ	�-��|Y$�-������JY�������	.� a.�I�Zi2��`�M� ���olKikS��MR�R ����?kKvI��li��v�8ɚ>����:|D���KL������7�R٤��y��의�����9N��u��%nO����g�V)u�S���ޫ�nݾ��~O-ޫ_"�=�iq��yUps��D
�����MumKK�Kk<,��}�p$X�	&\�."Y&�C���,#��x����ɍn3����;0x�,��	}\g|�W����K�^��%N���-�uq
94�w-c��1ϓ֐�x���x	b�f�-�]ޕy��c��1�A�����!'N���_z�lpy{�zX�A����A����S�x��A�3�P���Ҋt.vʨ
���,/n�\}�+��JvS�L����-�֟g��C̱=jL6v�v��g8�<��Y�>ɖiw�0��+�	��}��"�!���&xQ��R|̯�T�l��c��U��V��ڍ�r���eL]���Q�,��Ҏ
'0����@���BUUk��W-Ԩ�ܝ;d&
w��|M��;rzk��wt�����s����b���LN�K�~����;�~H�Q|HD 1\��z��$	�J�J��76$Ͼ��|��g��3�1VM�ܚ��7�W�01>A�[��]GQt����Jp�sK��m�q�>��ϑ��;���||႙K�8�)��X{X�z� |t�P��.������Fe��Ռ�|�t�}���X��A����Y��jbm�������]U#K[kI�W=��gVZjrr�|]-�ѣG�;��`�Q|G�mY��+�V����Pq�!������z,�R?��ږ��9&�������<�.k�[�glP�*١�=Y����V릩��H�'%V��k��&f��]�ᰃ�+�wn����J��L�>O������|����)�	$<&�W|����JQ
*`�?�NP�M��37e+�-w֖�?��~��
�6�YSa�j,�c�`G]]R�������T�(p7�r���5�8��2~\B�E{����������o�f��ҋ���@HЅܷ��F�oh�d��>�u�a��	Ru*ćê��������ShQ☝���}DB��fC�Ф�e�W�*���n�5h�f�Wd٩��D��,^d�8%ق�Y�ʃ.����Z��h����Skơ��Xj@�#6���ѽ9���Ϫuuw���Ǐ�G�1#�!��7�)n�Z�Q4�-i`n#&-i��*�Pr�	������_��.�~�M��Y�c��,�'�1q�И\��kCB"��m��򹂺'�l�oc�9>��5Բe�s��\G�V�1]��q{N���(8 ���3s�����qpA#�����k#�Q+�O���o^�����F�	������M�2�B$�����}>'ޤ ��4A�ܼ����ȐY2�@�����WW+Pk2K;�V�O}FN=�m���޻w�bt��iN�1�t���={�ك�v�?�1�n��}h�-��ظ�w@���Թ/�S��_	�M0'�D�� �#=!�Kt�4Lߟk��P��A)4c4�N�f���H�sk��iW$6q���6CD�+��DNW�WVc�D�`����iCF.��X���(m7�<�ģ�Q-��!$��+Cg)h���G��1�50��1�HD8�/潧[^�$�\�ҥ����!B��;;�PFF��ȵe���G���?���euew�wp��?9�-{4������%��Iq�+�F�/b\�����L&)��8|�tNv�B����8�uQD4����LP6�t3,�n�S��B���[K)i��(؉���D�Λ֏F�/���q�H�l��TH1g�%�A�	�,���}�y<X����Kp�s�kR7�Q�#�A�fX$�.�Y���Ķ�y՚�,��*�I��L.j\�фƟk��U	 � ��	���{Բ�p�.y���L�]��a����uS+��E�	ڽ�[2�js�f��\ē&���~�3�f�Y�g*�H|��E�g�F�HZ�>(�����;����xH-��=��s	��[�L�A���\]���i������^�r��2�N�"�<�lݤ�_������ܾF6v� !�]21�&�]*��n�oؚ�~��_���L�q1�5���Q��a��!�$�Q����H���-C)��0�a��q9��͆y��3��H����4�r����a<�[�[6h-�˸U��iG��Q��������ϫ����S��-f���r�'kv���yZ�+�vL4��r��X���Q������]ݷo?�53�g)���`z�s���+W�#?�Z�� �����8������˄��@l��:�D����ݰ��𓱪�v���g���f-��g?Υ��؎;����ɀ�}˺Ŝ֔0v9��קeiqA���Y��:"\aYF������FU`St�U�5�����_X��w�2���!W ���`:dyGMH&u:$]2t@ĥ.�6�Y��-�Z,S�Al��Xrhnf�B��+	��284"}]=��1He 1c������d�"�~%~��i��Q�b�Mf�A�KE�m��%���`H[�����B�݄A�S�	�1�p��6�I����j���g����K��׆���w�0���߫na׮�G�|qq����ށ^��H�� օ�qϞIV�U�'��F�?��h�ql�BW��9 '1���T*����X����+C�~���>;�I1���峴�8�� hl�簜�IT����>��lM3�@���2��7�Jm�^��(?d[�S<p?$\��Db�gG����$�� @�}�R�)H��`X�P~��h��=��1ۮ���#yO���N��n�Hpֿ�e=	J�)/���5(�-t�J�GQF��j�nu�����ڒ��e&6�A�J3VcQ�n�C�Z[4Uâ��X+�
ˑb��P�oE���Ji3Ȯc2pI�7��v~����f�Eu��dѸ+���a��͙�:�����}I-���g���vt}��<���$�� ��e\X�cd�m�?�A0�=D���Ȣ`�,�e�e��b.��}m��M7C��h���a,��ɗ|�Ũ��x6�'#�D�{ےs��;����ȉ�hp����ӷiS��0 �zO���ħ�%�@c�����@�@�'jC%��~X���ҡ�#�hag��e`���,/,�Ή�an߼�1�y
5p�X����(��r�-M!٧INeF)@Xk�=�Mv
�n��;ed�G.o�$� �ڰ��6�5ܭ��RZ�6Q�bmH1��5��CC5�5#���d�����Ҿ�������v�t�׊���9�~;�Z��rnr"a�%�a%�(�m���xQ7f	�=OlQJ��n�a�Qm�׈�t�� ��)����Eo�����׿/���O4k�8yR^��W���K��ٷ���I6��Yq��e�
L1ܥ@�����s(Q�SL��
�]�"r��&��E�\;ڭ�X�YJ�pא�h�b^��7��lЩ��
�z�b�0Z���ֳ�6��{������АLMM1��bLB�j��5��N�T����kv��ey��o�g��a�(�Iu9�1Z5t8������H�惈��X��)S`�q]Ô�Z���,Ǝ������ܯ�@��}��h��� ��#'C�C�l�v�,n٧6}`hhvߎ�Bsq��%���.u�|�t�Xl6C�L�|��(�;�/RB�bsc�h6)���ߣ�I �{�\A1����~ŭ�u~�͇Kr��%�p�
a�){dQ�,WJ2�gL^y�R�58���N u��\�Nԝlq=�EYx �3��tdÖ�8*�^�z
h��Y?J~��n�֚�Ѻ�k�u� <I�Ȋ�1�����{��Ίy���'�I�T3��R��]=�A�AZ-W줧��xW;�cOP��:�9#����}r��	�����A�TN��;�z5	�d%	�C�ܨ)�B:���;�טsA0"헚���9B����Q�� i���OzTp
zh0��p$F����~m5t�dj�Xt�I����� �[�����o���Lf`m@O@�|	4��@����T��ȋb�H�t7����V�/=�Aw�=7��	�F�\��B
�[h����\{ԍ�����Yc"nP�.(뎪�oݺI[$[
����o�����>����[��,��݈���z��ũ4]�hC��G�+��ƆʊL������v��F�����X�dĸ��^β�AkX�K�}���	�<
�J��%eB|!9�d >���
q��h�3č�J�cKjj� ��Q�(���*A:�Fg!n(ߠ5+e�>�n��w(E��U�I�l����z��#�s�f��ˈ�Ā�,k,��T�aq�gg�l��FS5�тfL��''�l.��{�1K�E��Y`2��+~g�,�f�¶�;���r�����u��2%������l�t�&N��59GBc���@��=۞��U�G3α&(Zg��fHݞ��{z`�!�k_����˂*��¼��O�O>!{��3�X�h�N��>ژT)1ٸ`v��CdX�M��&���A���z9-�	y�p�\j=c)�Q�����s�zb3�~{�.�t���]�a�J��:>��5\ӡ�\L
�e2�	7F���C�1��)Yd#��C1��P:ڲ27��N�q���y�"�M�����T��k��Fk�կ~�1�����\�z��A��-��
j�N�"bX�k��!>�yR�S�	�EV���I�d�����\��T�����P7��3)}�������b�(21������p;�+ s#!ݽ#D���5��?�Q�W�H6��N}-�o|Pr}��pgY�;e)	i�S2��744 U��zH,$\!Y���;��&rZ~КleଦS6p�T��\���f�A��:�܉z���6�v>��-��z��p��\�r�q�Y�4�O�����ej䈟�f"����L�unWˊI�f=r�m�n4<bJ���,��Y���a'Z%����{}hsqoݍt6�#�0B�0F�VoŠ���Z=:w�,��L���`K�qYHgl�1��VL�ʂ��؂`�Ӟ�	�駞�j�ܫ����0����2�bM߫�[ ^������D&I(e[2�{�J��k�flI��y�x?Ƀ����=<�d�HxlfM�i&�;��?^�muq�`z�Ϩ���h���`a#�
�2��'}^J��A��0�>��A��������qfe�3�0�=|���Tr�XL��� �.����E�=c���H��@_I0�[\\�E�^�W��1Y�����܈�HwRV�y���z��>�wR9,���D�����f8S�-�롡��&7W��Z.pND2���VF��^����Q�G�f�o񟞁�����v�b�V63.����DbE�R��*"̨�MV���T��x��9��w?g�:�sXz�{m0���^֣��D"	�+W.SȖ�H�'�<�<̪�usZ]�n�����Hs�;��@�^�"?�ɏd|l��G�z&�ekk]��kz�a���R��>��j�Ә��ف�݌Cw�Vsi�(�̇=�M�f��ǆ�jv��
�(EӸ�~���7��t����So-�D`�`cY�K��dA�Z��XHU��7ʹ"ESC��90��t�u2�T�K�,��!%2�����c���m���+����iSZ�}A� �@Y�����a65��P�0TuI&DnݸI:9�`̻�z�pp�9�ny������Y"Xwx�*�?b�u�|;�Ǟ�]�A�
�M��Oru�ƴ�(db�_�����>\w��s��y�T$h`wm���?-�s�� ˇA�33�"��X�
��U�|�
��C�� n�g�)�Э�g����n
�^f�eI>��<k�c�r�P17�l�{v�n0T�j\�dQ-_���W	�c21�<�O��s�l{��5I���ڡ&�(l�U�\�MD=�-��%}8Ӽ�M�dU���N�=�_Q�5�.�8.�����������PkPC/[��o5�R�J�� g�;���)���1SN͛O�ģ�6��I���sL]����}�#������LK�Mi=<u*��غ)&B�2��靨rX�_�kW����Cc���!�q�����Yv2������*�F��B� H,D��*���Ui�̂�LQ�v�ִ�˲��}�֌~ݖ5��C##t%K�L���fM� �_�覣�����h�kom���0e�:����j32^JY��8�%2��L3 �L6�!�-nOr\	K���{�tB��-H.�\L��@u$G��Ɉ6-��oP��Vp�Fh��;�H�g���}���9Ԥ�/`��Ɩ����䡇� ]��&�{���by44#>Mkh�"-���H?;s�Jwb�^�}�6�MO_RK�)�]G��OB��3X���̢�7�������4	|�A̧���j@-w��X����4ţ��ɐ���e}�M��ZsH�+vL.)2��H�f8�1C������/�*�?�n����䯿��|<?+yh{��N9&G�.���r��)YQK��wr��7%מ��>%�ǧ̡��!�z�ڴܺs�s�F{��/�$���We��G�y�I���?�o��-���&�/   �:���t�0�$��+�p_�xQ�.��s�����β� <'bW�E<�^Н�����VAlh����I��u�ڇr��duu����{P?�@�i�$8�xm�-"C�F��y²M�j|	��qu�Vle�X���D�E�����C&��֦�ŐD�qʐ�Ҳ���:�9E��ŧ( ������T2��L��37�ƋS����m���P$�E�AV� ��~��1�T:L���˗��QvH�0��l'e�����ꝍ0TZWo��C��C\7��I�O,���>P#S���	9��Yy�o�#<v|R�N���.Ȏ���P��l���o��z{i�=���kPѧo��IiEM�����e���j�ۛ$�LM�e����)�m&�	a+Mmh�36%������x�e�\�������I�L�A��������O�o���lk�U�ڑL�!�b]rTdۥW��k_xY���s|���S�¶|t�C���.3�K���?+���o�xg�$��z���__ڟ���S�bIC�swN�]�f ����?�)g�� �~��4���m./.ɞ�=<~"��^� ����¾����3:`٧T����7ސ�����@� ~�S�����X�[��L�=��*��	:@�سf�8�,���(ܱ�\���+Ā���؞�+`�P��ۆa���D`p����� �r��u�b7q�7o���ˌ��+��g��ř8'P��������2Ƹı��]���U��޻�~�u��F!�~ ��[do�fH� v� �t�Yp�@X�=M�u�C��g?{KL�y���WYZ[� �f��?�G�P�qn�����v���-�[��Re���4�����b�ъg�\d���opl(^��!��:^w��-��Kl;��ijc>k�����[ݶ~qV�ڐ���'�)._���	KU���r�s2��A#[y���~gV.��@5ˎ.@�lk�}���/Bk�
e��?"�|��w���d~Ux��-HB2�̬���xID�ZP5D�I[�B§��s�D���$�Vm[��9��;J:[9r�0�5���z��M Ŧ��m���X(u�X˃�����(��o��������ˆ�*7��k@�|��/��)uX�.=`�Ra�˸�jS_{7�$aq�.K
k��&����v��aw����L��v,hoz��Gڒ'��2�B�+����K�YaH��t&�V�H�A8po�7n����o㜞�/Cw�f|�x�'ԫ.��.?��G=e�
Y���`�+)�~��*��ҧ
��C��D�҃z�1���7~,�*x�Q[�F9z����a��^��M�̈́\�qK�v4�s��Y`BO����v��J<�A�L�`8I�t�,�!hkX�p��:�o]��R�mk8nJ�]P
�	���V�ū�U礴�-���ximcE:���6���D�(L"6������I�Շ��b�N*���4�33�̡ctSB�^^w歷��~=�Eu5:pP�D�7eX��e���4&̘��c0&i�By[���f�QOvjT����BƧ&�՗_�Bg<h!z:����Ve�#��4�<��Aɦy�w(�O��E�믿.��_��}�-HQ���g�&f�〛Q�!�~��T�oq��T�\�������-F.i"�Ue�1N 2ѩ��j<�����]�A�|���a����eY�JQP ��u��;�Zu��G���.y�*��>�����%�V��jnq�X�Rk�̝9��;��=�^@�K)�L�> $
/_�¤��������g>'�S��G?����ZjI˦*O K�: '�|D�Q��m�����v�2�Ӕ;��h��=-祡��� ���ED��xrO.�A���DZ� 6e��)i�C�(�f�f�&Ք�;��/4�oX7sMݘK.��N�������5h���ץ�(s�<�m�jY4���{Qݐ��z��9�d]�gmeM�u�4��δ���y���dM�����Ǥ2��W^�=��R*�䣫����KR�-j�h�M	g�C�PШ�1$3�4�(t6�T�����?_|�t�A�ڮހ#��ԍ`��,b5�=On���z�8C7�������_���P���.�d�댦�.�E}S��Fc�R���4D;yw��e�&�@���k�[�(������y�c�0�V��~R�1�n��-m���ƇU����w��ȵ`�r�|/hA�<ӫ�{`�*4
��%x}���e��^zI-�cjL:����@-�ZPL���/d�{�1fE������~��j��-�n�|���g>RpH?�D١�X>����zv5�ˁi��c�,�D�-�6�pLLe�~.4�W,qL_��Q�)P��lZ�,���X���U�֍i����emaQ�����V5�̴�T{�X�^-����39��{u�𳪺"gμ'��y_V�5�
6���y۪� T���i�v��w%����z�J9�/:��L�%,�Pl�L����Tb�ժ!��^ِ��Ւ���~Z
%Ce״�]$�Y��POsƹog�����k��7��?ȝ�;������rl���!Lp��.��Ͻ�<*�����T�������09�;N�#�;P�T:���r�����haNc����R=����kZ���5���р�ͰXO�^pϠ�W� �?��.)�?����ʹs2%ђ*Md@O�>�f��x�_�ş�;?[]�uf���e9z|JN?���z�\�9��FH�8��.˛����o���6X
kh,����{8f���
�b0�����G�xgGYq0E�v�����ŗ�76�<�%��b�%n�^�%��,L���f,�4�zP�m��)�di~N��9���8�����.0⋵�5Ɂ��3ϩJj�1T�k���hSX?����Ե��k�vͪ[�.�?��?�}泟!�@,R/X��n3"��A����?�?��?�s�7� Sfv:��֬E��:�q��l���I$Y𞖋�Bs;]�i�Xԇ2XZSQ۴��1���au�8 ����w��[�k�R� G��[n>/��e�v��~bM�5w�(�νw%XĪm9��3�"s��߷o�0Q��/���ο���z�X\�lĂ�RG[��+W/ɟ�ٟ��o�C���p���d��y��r��^ΆD]���������9|�z/a��� �����8ˎ�Nr�,L���Ÿ,		�1g	``��� ��şM�ph���7�d����Z��K,P6���AM�w}�ބ44�<�5;�}bH胁�% D���u�!D�?��^u]�:Ĺ����e�z`0ݴaIh�uMÑ��b�?c�혩�&DJ}G7�P_Ω���������o~]��[_�+��iW��;i(��L����'�w�w��	k���~#h!r�L�@�#y%�"0X��L����t(�%�M���lDX�ڑd�{���Y��� @��Z�]g���9�[�Z,d3�+�d��;�� ��pJ�n��f2��z�
�q������^ܒ�C衤v�� ���-뙽=;+���Y~�����_$ґCU�r�۷n������|�[L� ����&c�C�9p`J-�q��P��2C�����'��hnV��s�Uݟm��U����6�IN��M�����Lt)����J?��6(ֽ�Q����EHS�PC����˘�Z�J��ҀsQc&RV0M�O9�3�`
"B�V,����r�X
A��l&�(,C۩��!�)
:V���%�R�P������5<0|���`�������?���=��9qB�����E�z�*�o�?���8�;�BT�+��w��|M����H�.���ErH'��˳
7����	���A��#����>�>�[ds��쮓�3+�`u�s�������w[����=�[��{��!�o:l�5`?��W��/����lcPJP2�6T)�e�vU�@t�?��c�t� +Ҁ��Gfv����MYV����$Da}�,xJzH+v.	�}4@'[f���DfW�/��~��B��ME-	��B���?����JLw�1��b^
k;j���)��kpU�`��k��`cS&A��DS��к!`�O��:6� �2o�9YB�s�x�6CǶ(O��$E<�V��?����`���Ɍ�ݚ���s��6�o�ؔ��j�wt��;F�/�>+��[�O��9�
��!]��6ƫ��Y\bt�c��<v��Kږi���:�,�}.
�ZI��@�x������}�}�V�S2����" ���k6LBgqz�^��vd9����������џ�cG����S}xN�]� U����[f�7䂺�0)�C�ܨJ	Ě�D`3��y��� ���"iqf
����L�O 2\��v�F�q3t�Mw�k�l=�'����p$�}��>s�i9�wc�55��k�<���V7h�n]��q��I��\�9�}�-�!�/�"1���i��z P���sry榀����9*�S�����;E��>�sC޻y��l�1B��Q�i�ҽ��=���-ٹS���ʉ�?#��YW,�mq>�m,��F=~`ag��?s�lnmp��χ% ��ۅ�l	������$ڄ�{����adT�~"^3.x$����E�t��ia3����?�Ȇs<��'�EmeFq.���+��h�r_K�8E\�|����e���f�"�������)�_���?D����^ɶe؊��Vm���2�� ͑ivf����V�GRmҝj���B�U�O"k���4�9M��dk[	�c�d-b���O���QЮW+&3��@�SV��D3�[f��;d�X_�6jI �}��/���������rA�U[ A���K~uY�DZ�}H��7�!��ݭ3#x��5�����r��U���������ߔ�jx����������d�V���!��/�*��׾!i=�;jqa���3�ӷ�)��oK-�Qsc�!�J�Y�AF5�v� h���Y�����[r`hL~��� ��h� ���a}s��z�t����s�Ow
 SM+��=*�@� h  �A� ����"����`bq��h�r��̑f�aN�.eb�] ��FQe�fa[H�4H��[�"3k�u�Y�\Wx����J�\G��L%���q��Hܽt��ڭ�����:$��o���b�(�z��a�lR�U��/S{������6v�����%Yښ��ֳ���Hj���v&!K�m��4#[j93�����5��%]52�#&̼#x�>"�$�L�Ag�o(P,nS�lBorku�Y�Ռ��H�1${���\w_H�	3u�T������PSߩZveq���Z۶�N�U����/��u]�v�'�v�46LK�� @_�5-�7�E|���:���ܼj��
OIR������خˇ���S��Cd]�Z�� �H���U��Q�"�B_�gطKA]
��PA�9;#��A��]2��׭�d��~v}l�oJ�Ʈ���36E�X���C�i�]�9��P�ͤk�؀��!�m�v9�����Lw0c,�v�؟ȹ����֋�jh&��V�.�c'=�`�C�<5Pfx� l�D�Ճ�u�Wk>_�5K��H�`ف�a�z�=~�E�/d5���S'TQ�ez�,�\'��"�
1�K��C=���n���JYyU0�p���e�.T�[�GVQ�0L1�}Ƅ.R�0��r��|1�F��>���#�\�����Y�X7�91nF�{p����sN3�exrB�=|LΝ=��nC�:*�\v�
�����;����O<!�*4�FN�_���?�xF��LR�z���Zn鄺z�m� {�}�GZ�>}�#�l�YY"��S��ŋ����z�1c.���u��9��;����򙄩��Ar�^�|#/k�B�5U�6i]�J]:�������чeD]�����d{cc�H�h+l���W(��p29<�jyd}˘e2�q7��á���+hܮ&S�΂��Y��oc�Ac4�S"1�w������F��09̰��������H�C�5��1/c��0�JP��g��qJ���"�sؽS{���=�#r��3�N.j�)��n��jRlT��)-�I]�*lx$�m�)ܗ.}�v�p��R�Ph���b��a?j����f��Ĵb������t$��"0ZZ�3x�tBR>%�}8S�}��{�5�2:<B�ݙ�M�G���3�>�'M��>xO.M_�������2�A0|�2�L<�ß�zI������,��jQn�.�P�$��mF}�?���� �3p�u�c�W�e�����IW�r�V���f�WH��%k�j'�96���$��冺���E�T��t��5�����Ĥx����K��*��S-��8��i��]|v<��&�1#^��uY����j���b���O$|H��U���c[P{��ͭu���w;� 4�����im=���V��c�m�y#��+�Z�N&��a�P&�,s7Ja��q/<��X;��@#�5��W�ר�˝mrckUT�)�Pt�8Y���z� IH�h�0+��rP�$02�;\�����6��N�uY�]zF
�h��]��7m*D����ݭ�K��̜�Ǵ�A��`WKM��i2�����(��0ɨ����,Cl��E��x�E��+�:nmm��ڒZ��k�)���Y9����dA2_�p�A�ڐ�҆�,�a�F�W� 
����#��f4@�Z��Z���>u?�ƅ@vL�7�#]�R]��0.
��A��A�����������u�z:$�q}�=�{�⍙oN�9�^+�\+*�ܰ���O6*7L6�L���*��z������@�`�`���U�=��:s�J!邮RR�l�q}��wc�<�DҌK,�͹��F���qa�[� &̻��������@ל�K�cZ����D���)�.U����5&�:���5ܳz+]�Ƈ����ec�"�K�j�����R^D��ӣ������G��G��-58%�`�n�ǖ��>�ɇn��E7>eF=C���f��'d;=;��kQ��ݬ�es3���k�H�<LAH��'/�ץ<]���&NIȁ��hF�Pέ,���Ac��6d�+����	�8�ԵM�	�,8����\�	�,a��v��76qU]F=xzO bJ�����J3h�k�+x�F9/s��-��^�T���E�^����E>އ�#Zn>b3CLd��}R���d"0�r¶��:>8��fU���Wޒ;}Z��L]����l�	,��= �p����8��������n`H�{�����0�K��%|*��z2R��d]=���%�JC�u��Sa��t;r��!y�cr��U�n��8�q��Կ/zr��,-�a��^�l���ru{U H���d�I�.&4��A"pA���[7I��JL� ��b��Z?f�|�4M��]� �h�2*�d�
�k��$s>ߛm-��d�Tb�*�i�&�PA���(e�"��$9
�����P���4��l�t>��,Vhռ\�4c:Tt�7K5� @1����ߴ����(���ؐr~P4#s\���^SK�/� v�:�؎�A;6�J<��)�M� �Ê�&N��=аj!�Ϲ\�����xH��f�K[b������}p�04���q�9��
>I��uq6��tu��ΠS.�Q@�I@��|�,;ۖ�l9Й�%Q)�nN�Q���n9qdBz�)V��g�_�y�����Z�b~S�,�+A5�g�K�8yH:��U���RCz���*nK1i¤d��r��sy�k��#蓈�֚��j��#������'q0Q�&a�m9"4�����$�ί�9�t��V�"�1T{��:;u1�p��>��~M�dǃ��_M����r�T@B;��<�L�Q�;�%�_�ƨ�*�P���!�X_i�p�'�w:��֎�wwI��S��
c�v2T�U[���3|�n��0�}��@HQc[�.�n�:?��)~��h���*�h\px<v���tS�����}�-Z�"x9}ʏxIq%lg\[71	n*�(�	B�. �{zzٱ�5�\|�Qf	����''u◛OH��5vYU����HN�dj�èi���*hU�~��~A����<�L���I�t{~NV�_���˩�A��2��%�� ���*+_��P-�ճ���W�4V�B3��ѯִ�C���[+F7�M	 ܄�1\24@W>��Ű>4IC��	@+d�s#�_C.p�N	M1���*��}��u��S����V��&a� ��.C�R2�h�&�/j�q����iS����i����ig���A�uu�?w�����{�./KV��/���t��`�T+.��D���+�7���|��Ix�'fι��Zм�ω����KC�д0��[0X�@�LVRl��,r�le�b�f� |f��4�#�qh7�d>���#��\?�����d��XR1�+�uZ}ux- e���<���d��Lq�U�@h����).䁅��>���1�|r4lQ����iY�V��D�i��E�1&5��4���(r_��M���=�rd�W�Ϯ�Fg�GV�ԅ��/�\��4��6sM6*y5}\(�UD�~V(:�L=ziISLpIsP�˅<6��MC�ql-(�֟���&~E��K{���,)0�=Ã��;I;6q��F��_u?g �
�9�Zݸ����Z��Jy�T`�AΑ���#w%x"+�`���DS�7�͆�C@���^h����@�#SYGIrzh���{Hzdr�1}�W�Z�,��	#�"
�8A�Z�&c8���g�dp���tt��g���u��&(�,i5ɊR�h������(���fl|鄘DKn��~O�@<�kAۀ�ad2>�l'�z�<<x��#4��@�x~�3r����O6QM.c�b�Z^<9"vv*�랡�n=b��) <��cS/�����RC�$,#��� �4ӹ����߾0-W��e�dH�ڳmr��<�.��N9��)Y>��}�����٬H=��K�i]�h�y�f��[3w=e�$����ψ�|3���Q�?\��ʆ���FpЮx��Լc�:{�eysM-�R/�Q_ Go��!)���]-��w����e̽C�����]<�� e(�	��7IS�x�sҹ¦)�J)a�#0]��Z�١� ��:����,�7(�(ЦQS7�>b>]j�)-�ܩf�f�6'��!G�w�$,��&m���t���sZ�<�J���g�s�{�4�w���GK��!���ơ�m����0�$Za$�)۫�L�7!i�1�lt2ؙz..sP�,g�7�B0�h�U���+�kź_hz���G�#�Yt�[Ì�ȹ�==L45�%NU��c�1y�Q�tM�/#�ɪ
���yY�|�T�$b�.o����O?$C�ސ�*��>+r����Ꞵ��TA�~H%# 5c��9���.K��KX���p3Q �l�:��b���4��4��&"ҾI7��f�wqc[�W�hM�{Z�����E]5�@��5�H��ɪ�9�ܮ��Zg��ʊ����
yʶ��BӎԴ�,��<G��V94�Q@t��1l�5&T�| ��P�7��{h�\��膉uC��2��J����.Z���n�Z\���ũɨ����%�Q��2}���P0e`S���:{x q�;Z8˹�Ho�1u)�O��H�6-6�Ɔ`�[��k㉻{%����N�D>�Q?�>l5K��A�:D�Xk�xF��qYR&R�k��~�%Wc�_h�B���)��z���5���F�"���������r�Ί���������}�|���J������$�=�%��`e�����uI	
�-��X��l��/M��d�Bl�2�&�}DU'C��4S�J����G7G���U
;
���#_3��`�LfE�th�Bt�v�RhS��,	tI-I!�Z��
h�&m�hl���/�Yph���	��b溋��`ݐ(��1B���U]�R� �ǎ����!N���B6#���<^@�
l	���B��<���]�8����& R �p6��;" Z�&��Y��Z,��ƥ�DB�gc������ZTr�#�,���N��j3mPQ�8�o
>DMU� |���9�ܚu��$�;ji���_��ġ2�K�YȦ��s�oz��ι�XO7��	��ַn:f�����B�Y��WҧW�V����d~��!~*Ꞅm*6vyr���%L/ZlTevcK�a���=2����}Y�4�m����M���,�vH���Bt�C�5��g'u>��ll��q
����?�?%,#�A��E^��<Mv�C�f���(?`$W�1�~͐K4��ɨ���ZZzfn�I�l�]-c��&E�2#{����3G�k�8)a�6Mg �(�m�<�.�O�����o�7���o�`��
�G$���w�����Y�sE`(3ğ�D�@m���y�mդO�����T�x.��h|���X���=��V&m��Hz����'�
��}�_��5.�B�fμ�X�r �����6̜6�%��\�ctn}���A�PO�t��*�|�����ӊE�|�f�>4�/gU�A45�]�GAi�Pd��/OFu�`O�>7n�J���Y���9�Kg>��|��~���IQ?�K���\����i��%]�����)�U07{r�ڙ�j/�q f�kd�l9�k�?����;l���Y,��Rp�<�O4)�`���4��Gg'J�kD�f��@��C7�`�%Hl�R�Xc��Մz͚�;%���P���eim]�aE¶-��Ԇv������Z�-�{�P.�N	�S���C�ıG���E��U����l{�L��=���o���|�����'�N.ݚ��G%��񺰐���";U������f��N/�t}��x��0e�&�0� c�G�Gغ�o�~2i��
-L�t�����w����)B`р��"�}�B����$bV#��lN�I8DƱn�;5%��{�����̐����qH]\��͏��/<�
���/��#��\i�?�i�rP�)�����P �3�+b�R�Q��M�u9s�Z򲺶�N=����������W�s^�dG�Żf��ś�-6(^6'�ȓt�H3��luҔ��\<
I�o�xa����4�hϴ��_���������b&��Ѐ��H*���RX\|h|�`[���nL���*ku��q��P�@�f5�Ù�I]z��H���MF03���t2GO��8>l<y3��.4����k>��g����'�}�2{�
I{s�)�{��M�`O�����"���Gr~�2A�Pph�4�$�8��/ļ��k\K�C�.�o:�[��=���t}��Qy�����C&iPop^�(��m�C�����	�{<���d	���s���̍C;;�և`8떱�1G�D�h>���pn�P���h������-��� �
�&�2��I��A7�ݕ5���L�WU�Q*�Z!/�z�#I�A�*;��P�QOK���G���o�_yE�rR��ܗ�͟�B���+�p�:��E��/�>��������|���'igrs�TP�z��ά�}z�F��}˗~R�#��������*_���~u��v�`1�!^�.n�Lvz���������M٪���a(�60��u+äo�����U�$;�g$M�I�Ni�6�l��swcH~ e��Iך���^��Ka}S�፟�����KZ��H�Kw_�<w�i�Zݐks���L�`fz�����15_]t�ooS���ҖS�
b��Ȕ�LLߞ+����d�(׭�J�!-FG�/����ő῰.�%�0X���,ٜq�!���A` t.�,!,#\]w���B�jB���R��|��B�r;ǁ57����B�6���!
����� �X�g� b��y3=�)6dP��N�U�����R/jJe#�o$���)z�r~��i���ɓ�:&Sc#�P�4��d����Ԥ�~[�|�R������^�gW��b�zm�'0�	��(#`xt�d�9��������u9*�ңo��'�~�����e׿�6�i���y~Z:%ԯ�s�>)o���|��ʭ�;���0����-;�*s,���IƠA�0r��a��NȬ��]�/~����ڥNËO~V�y�Q��kߔ���8�,�zO?zJ���a�f�/^b�:FG�w���ʋ�{V���cuA=����/��{�²���ZQuG�1�gʏ�i��rڴ�d��,��1�R�e��4� �\����*r��{���C��{���R��_�n:D,^4��{�t(�U4s8L�?#�������E{���'�p� ��o�< �K.�\�L�m��>}����w����"��d��#��������g�<)}݃Ү1���y��Q�?���� *�56,�3�O�P_���x^��W������	Uf�0�Y�V#���!��m B�I�H��)��z\��c/�#*x�N�3j r��?���V���ZM���&"�.�W���L��׾���_�c4�>pJ-�e�z4h�a�
����b���E�H�_��D)����Qm67s[�\� �-_|�yy����ϦV��y='y�i����z��1<>*C�ҵ� ���1K!mxDC�F �7�ͯ���"�
6��n�/[j�Q�Z����<L�A�${C�XK�����2�nmu�t�g3���|����{�f��j3ѭCn�8x�\,H j��ja�X�@�.o��$�M��������~�"��B|
%���$��&G�ՒvV�VEّ��NN쑧{\�= ���9x��׸}yy�Vwep��)����oW���g��7~D����!:X�3�=釭��vIK���Hi@9 �����\��G%N�T��Y��"�rW����]�-G4�ek�L��[^F�wL�~�_5J���G?��j$�IjoIT���ݜKθ����'��U,���Cv�M-Өj���eY^���<�|�!Ga�)��;XG2X���A����λ��;�+}]294*��[j�(�T�qmR��W��T��n��a����ls�ϰ��ZYqHX!2V[�YNJY7��A4n�,�xLڸyQ�m;A4jB��j��%j�["g� 0�~o#re&�l�4^�+Z�� ��b���I��
���7k�1{�*����=)�	!�%���d�*�gB�����<q��=h��-��ʕt��Pw8�����_=�����}��/�ɓ��;?����w�I����e�#rH�6����*8A�<�S�B�OJW��Z���r��]�:��8u�}���)��i�1�c�;@>50*_�̋�����ے_�E
��6Y&f��u_�z�a2���|����Bgޟ���o�x�g}m�솟�ܒ�'O�7��59���e~aQ���#���:-��O�{��v��7�)Ս<')U���.x��ri�}�����a��?�8j�!��ġ�ժ�A�\��L�X[�'��>k�RF� �~ps��	�C�`ո{T
V�����B"��,��1Ŷ)�=6��Nx���1���	!\U/�/lm�k�����dv�b��%A?����Z��Q>�z![�����J�sRN�>!������@� ;k><wV��ehtD*�
��`���wb�O=.�zY:�{���[���_�Nu���{�Mn&�h�9	9�Z�<���#|Sly�P�%L�<K�+_�F�p���ߤ<�����Ɗ�f��7�R2�
�rz���͋���}�Ţ����K�/ok�H�~��S�;�� �W�J]T��.���t�
�^�.�#�zN��Փ>������Y�v銤���p��4���ٙ�j������]���>}Ï1P��.~JW$w)ub%�7oh&�_�:��u���ɶ|)$�h�:L��G�����2޻�y��i����0I�Т�⍼q6n-� ��n�A���a��R�ߣ�� ��r��gg���oor
U	�\�3�|����WƆGd�ظ��j���q����N>|B���?���nʝ�9Z?<��zI����SOʣꪶ������~F���|�ڻR�.� 6$Y!i����ne݌�ZQ4�d����_mp�=[.w�)Z�mM����g���}����crsu��p�@�n�L��A�{_�h�lm.)����[/U��Q������N?��@��+
N�w�{O~q�}���`�QgF���ƨ����dz���(3����o� ]� mm�[���!����C�|�r��/�A`Kz��-�.��t�?ÉRi�-�Xv@M�~W�d��Ѣ�V�&�nϺNG[�w�]���8��u�i$(�U	����}�efj�*'�',S�ˇ�Gf�5
���>>���L�����y���O�=��I+%���j����W�Z�ѱ	B֮^�¬<���.k��eE=�����U
��_z�U�O���G�f�]��-pg��a�%_ޔ�[��vcU:���d=�M��d3���v��=����H���U[)��T:�3r��A9{��l�W��!9M`Hq�_�2�8/�o�b>�nJ�T�"�c���CIow��-/�F�ͽ�����	��*ǀ������7hq����HwW���'T���#�}��W�J9��F�<�>�r)֎<�v��sp���il�h�0�.[�',�Y+B����L�1q�ZX�Z���"Zf0�ʡ�<:���̾�D�2����$���ۑ�����l>k��=�~��!��`A%��D��[^_��RA���4<��OP(�D�|�ǎ���1Z$��L�>�d�j5�ߚ�۳3���N��?ʡ�j9!OH�a䷟�Ho�C�O����d��`:�IW�ن"b����e��*?�m�?�݇^�#�/9�l��'����k	Tkӝ@��fXc� ��͈ ���ew����')�����=��r��_� �s�`B��"���F|�b�%*`Ϣo-��!jd"A7 <2'O?*S���9Q��#fw���9}M6f֥ȩ5�~q�D�d��$�����OJ��;��j%�z����d�2���V�qN�~Iv/�ea��V�����$����[���]��>�J����4��$\܊��,bx%��C��B���c:��bȖ���=�[#��8�n��	Un��S>��ֽ��T��FX_���d�f;(�A��1L򅒞�Z���*[�h��i�N�6,llI
�wP�G��--���X[Q�$'�����)�N�Яi~��)9���GF4�K1LY ���Y�[9�o��8"�*K��l'I��4jl�E�tѫ��/�M�W�>-�:ƥ�o'}��ݮ�y+3*%�b��L�)2�^���s�S�h��TT�p�Ғ�'e�i��Q�]2��G>�&��7�k�l�5��R?,jm�BY݅qy��g婧�"�^�Rl�K��$Cj?L˪����vTZ'�V�Z��)9]x����F�[#���ƌ������*��nh,�c�y����;�"ѡk�QP8v�tڡ��NrqE�v�P���k1rM�.�s���d{�ȸ��;�\�{hC��sU�0�MҎgBq����o�"�yf�9 �k5rn�|��u_eS)�� �Jg5X���؂��kW+����6��Os6����0��a"1&c�د��W	 \C�^^t�:4�@smn)٢43��æ\i2�L%���n�HΝ�(�F&��I��;�鎴0�_�h6���h`]c/�Hw�C�;*�O�����}���q�H��!}�^4,6U�=kܜ3{��t_Gw�k�Ќ��𤻷[T��U�|}��nh&������;"j ?	H���u�������S255%{9�����+�Z���^b�vP(��'��,�4s���X�]d������2��)5�J���Ϙ"7[��~��c��hM�����q��-h��?3�yg�+N��
�[�:��z�؍���ص�Q�&v�;j��uF��%��H�b2�!CŲ�ðU����39
P+��Uk�XN��9_l������f0f7��8*��#����e�SO��쾈:�-���W�O��F��Òe=�9]���wdu�*G�6z�aL��X�f�F8�4� ,k�ildW�Sn.βg����vI+�w���>��!�aѺ@�Y� �j��s1��. 3ju��>`fv1
���V+8J�\� �4jmm�Y5T��x��W��3.�H��.�.UA��dCݝJ�D�v�ƌp[���(��$:,B� T踠��a�	vv'�Y8p@���2�>[������c	���f2��y���i=�(��4L�s[�?���q�N&��k�U3�f�\��~����'�����_G�Kh�Q]�
�V67�sB�@ݧ,��7�C�6�"�>@H�t�HF�.���>����^#�}��h<YR�O�4��,���%�RI6*5)�lz��Svr���M}���B�SݍlR�i�A"�V��J
�"��b�9\84�|�!��%�Oe]U���z�Q>޾#�X�*G&H�W�`����l�b��Z���e����[�����f^�i^}��b��� �������6ء�iT�r��O�<�s�){T����	��� �����h��*��FxS]ǭ�u*�����L��C�O��}zxQ����"�0-e(N�E�?>o/4�H��F�6CTd�Y�O�Y�zJ?'�����#�<��G�nK̭�t=t8W�Z9z���'^�w��(��k)*�uw/_덌��P1��RD²VO_��sR+V����!���uzcsK���9�����nl��uI�X��ͼ���w
%<��
��XP@Ͷ�=�r�V��+�Л�.--q�Ud����L�L#dshm1/��Y���x��Ro��<�x���l~��ob����P�,?��=���|���O�.�aEfk�Zٔ��v���fS���Ft�u	�� �`�Lq����V���>��r�:_"��e�T��4p��d���R�%,��0�KzueY677��*ĂH�#Y�hH����d��Mӏ�_�P��jK�go��1�Ԗm��z�x��5��-���fH���!�-��c��x�rP疁�ϔ!�b��=Ɍkz�@84�&�;�fY��=���odUc1ۯr�F�&;L�:��i���5I(�űw/�{Z3S~���j,�3[F�"����5j*ly�_X�B�.>_�Z�w�~G�^��!à��c����}7�����0����!�fmk���^�=BjF�K�o��[ipv\�;-�PD��I=�.�Х	C��?�����oׇ��'�-��i���9�f�AM�eecE�Ǧ$�%"؛������
B�L��c�� `���`���u�u3�u ������=: ȅKҨҲaQ�|�کԍ%���`+����Y�2=�÷g��9y����J�����'���^3^��b��a�*�:&Bե�W�C���o\sz��e����Ic].˵��׈���%
��;;)@(�8O �+M8K�,qF������ Hw�q�s��Ok�B/����I�ΊF�-�?�5�� �Scm H�	�	Ө` ����y�6�ܑ%�2�g�|��ŋe;_ �Wo��k���ߐ7�}�'�����5��5O6v6�����L����҇K�˓���bE:{�w�C�Ќt������57��� s��aN�ۨ�"b�Qm���D2	h遢~�4M� ���L��`a +���>#�'dH#� ���ˀ���?��+J�����#R���Z��	�	$Hv�l�����ؿ���ܿٿ�=�{�Lo���f�lJ�h�кP@i��R��:�׮����"�3g��X����gf�̮]�.fp��
9%��(�2z���ƍ��(��EM�zޮz6�۰�س��(�����6�*�`�0���oh��Սl!�3k�/-��u�pG�T��f����j` G���#K~�&����:QZLɢ#��Rrd�UXX�Gna@|nϝ(�v��܉?��6'
xH��m2��[���9���yP�`gP$��8�أ+��MM��d����t�x�vG��_*MARt�XR��-bGt@qRڪ5���H�� �o�\�d~��e,�,b�`�8+1@I�z��`p�&��38s�.]���v�<�7���cX��a�fni�������#�m}�(ESDv$��,���N/��fX׽	�le�4��Mr�g����U��r�.�U~�iE<х�t�����^�Q��u1"����P��o�C�D�z�8Y1���"�p�޹���OrS�a�x̨f��]�����@fBŁ�~�d�W�]�jk�V1S��c[=#��0yW�-��+��5~����Ճ����nؼ	�7�MOL⮻�B�@ǥ�E;�VQ���׮b�ƘF�ls�Y\��ۋ�����k���J���i��MqSfUiZ�J��C�����V6ͪm�J�TgՌ+� 2;V^��P��ۭ?�L���v#�W;�k��jS�~�� �k/��A��Wm��f�ANd5�:hq΅_Z�D��\WP���OLNb�<3EO�'1'�g �ݩ���;6jFa 3��O?��=�D�,�̣P]��������kN�9��2R�R���,�P���}@�(\�9>u��c�묡�R*�k$�L��#q��ۄ.Y�tCU1P�	]�!��(�J	?v�z}V�B�DE��M���$<��w�>98�Q�U�K8�#�ԑ��ЮC�w�+܉�����)�w������E������Գn'!9SRw�H$�(CƂ�x���l��5uy���7���)e+r����ׯ�̅��/9;5�?�ۣ^KR^�p'���#�҂��m�5��S�5��OMbY"����X̬H�W׹Ee���)�/U�3ƑlHnVm(�^�k���a�����;��Ѫ{��n��}K�ir#۞�I���U���NS�����g �ڍTWV[����`��~���H���A;!Q���a��]t^��J��ͅ�[�������)t�	\G�ٷ:���WPϧ��c����C����-;�G?'�~�z��������
��d��naI�	�����˧q����.qj��\����УV�֗E�:�!��f3�<�0Ώ�#��,�+��E�v�
p��qeT[?��Oe�c>"�z�&Ik�E�r#ϔ'qc�_����0,���Keǯ��bnyI7�R"���c߆-�p[mF~�,���r��3��qێ]�9��܂8�%���P�5d4H�8ka%��K璕w?��v�@UlR���u�Pr-y$ޮ��]�P��o�g�r�3ٌ$�+�[x�]������:5E	T ��MB�~݄S�(�W	��0죀����-XP��oU�^��96�Ԃ�Yn���\mT[=�d�uۿh<��Y�����v��r|s���~�u@x�BGC6���|i$�ל����WR�Ay>+���|Z"9�a����'������Ǟ��I�:�:<]�gu#�g�*(GH)�B��1��DA�Uqt9a�~I3�z�ju�7Z��fC��'1$�aeq=Q����zB��<��̈́ʦ-ai=Ou�V�TSu�
�uJ�塞B\n�@01j�Η�r���>=i6�z����d���doڍW��4>x�8z�~���8?5��D��֋�=t�=�o�AH���x���x��ǘ�,!֓B=�2��U3������(�>�#�v�f��%��V�Yw����;�]AsY��KjP	X)�$��(��C�D��l2�r/Bc����e���j��v5*bvć�Ls3˹�◃Ռ����vl���m���7�e~S�m�ʩ��y~�+����"��o9��`_�VT��w�L�"�Z�}����QS�S�܄�➌*��G*��+țYLc�K���¬8�E�`��lE��OE%z��Z���/O#$�i��-X��e�̈���(Ρ��O
.�O�J�KNW� ����bA�fy�ID�Q-�P#4����p���J�#o��λ�7]����26���n]*ª`z9����G�ͭ���l5���T��b/o�/Џ���i��k�߱��Y^gAǫ��B�5�k48S�����Ɓ5��c�³���|:�G�} �����~�+�����p������#O
��N&�ݷ܆=��G��e�>9���BuV+��0+����Gq��=زE���E,�/�v��I���¶W�M9��ڋ�����fWT���tΉ�IއU��$�Q#�07;+�⒙@���i���Ϛ#��\�H���h��[��l6�=K�����@��V����e�g�:/�ڀn�U�!}ߚ�΄�d�F�V�E3_&(�Er���you��<�����{Ͻ���Ou=9�$��0=�㒮�p��ILKηn�Z�`g&t9,�uY`�+F�b����I����2��gN)��m��bߔ��j��P�~��O� ����]��ؾ	��&��ӃZ����t� �.��0�����W�ZV�Xʽ�ꛢ���1<uߣx�߿��}�~~�}]��w`��M�><��c�!|`�r0g�0/ƿ�� ¥�*|�X�RU^^͞���ch�ʯm�k�}C�JU��
�;.�;tX��"~��k��#򬚴ǆ��gF>˙+����}�f��،EI�s+�[�%r)3�zj_�	9�D� a'7�:�la�ڡ\0�����R	���
�&'�(G�F8h�{ڛέ����n\F��%2Pɘ�U6Gſ�u3�������V�Uߧ��i���|D��X�9��������I�݄��4���l������ºY��H7:7�E��#3SJkL&;�ܿ���d2��ݨ�H{�+�ke���jT-Kr��������e1<?,�+簚[�p|��.`fqJ��nW����FHb�uM�k8�hR�sL;�G�/C�v�1�-J^4��DU�:��D���><������"��!Q��Kcx���x���a5U�y�I��4��h����������Ѷ�A�$�,������6�F�	���i��8����
����Dy�TJg��./����u�M�@'e�{$_�7Z�i��lx:��/zCzG�8�+,���Ǳ��r�qX���%���y�`G�L	��
	�q�쓵}���;�[���b���P��N�Nz�әQpHBm;�����Z��0���n���^�U"WCl|}86`��1�5_��V_Dl��FM���f�{�M;��G� C�B �5�=�e��L���SUwmH4� PtW��������QGE�����;�����ae��J^�,�mvi
˅��a$:��	�^I�t�nmi7Xvo���Y�i�Q|[j���fk�p��	���%V$D��x|IH���s���fݘ�I�bs�{���#�%��=rS&/_��P
w�ڧ����w
N��۟}�1q����կ������>��DJ�:����i|u�8榦�3c_$���j�$�^,��͚w��ΕsX�����z�Q�)_�i�ƞOXǒ̬᧟��و[X�fE-�ug_�Z��*��8��P'E�1�����i�{�XA*ߊ ���[��XN����+�Ѷ����U �i�� �`/68��f�0|u*�t��1 EЏ�?�ᢑ/�6��A��V�w��t��k#A@H����A�Z��n�D/2��+�hhC5l}�A�^�:!��yJ��d��MӺ��r�r~\	�o��/�*��A�-; *�ǹ�PGq�@g���H:��nE"E��������Q�@yҰ�J�gg����[Z~�*��y���!��̏XZ��֋f���b����%8��=���^[w� ���)L��@9� g`B�Z�6&p��F"���$F�_V�������ȥs�$8���������E�}N��i�R�>���M�+1��-�m�l��>���9NXЦ�Pn�����e0�6�L���+a!SB,ihf�<��	��j��YP�z-6��CX	�E�-�e�]4l�%�/��� ���R(�{��C������4,��$EP�w�9Z�7�y��Su#��a1�eSڵB�f�*6��lku�3d�`v��kUd)�Lcj
C��ߨ�*��_N����X���`?[���Ir]B$.N�CΨ�7���R\C,���u��\��I���$�.a�p���S�4��t�#�[�ԃ|#_W�U�|��+�*�rt �\�Y��:Gp��Ɩ۰i� �u�˳�� "Q�Qk`ӆ���w��f�,��ė_���?���˸16�zfq9D��9dgg��с�8�Y���A�ULJ�v��9���CMr7:�5�6�:#��vj�
�������N~�Jih�?��$#�@i�Y%S�f��%�:!��<��|�:�ȗ�s�^�ݱ�׮����X��9@��vۆo���f@sL��a#��nsa�eh~���t4����5]�e�o�=��-h�a�Q�UEuVg��K7�*�gVcM9�A��NYHt�e9KF�(d�n忾Maڿ�݀c V����;�a	
f�%��A�{�f��1�,���=��B[��rO�8���q�3�i�f�k]������X��ȴ���������b�q'��p!����@�����I�[	�ٮm=� 
�'��!�� �����w��_p������.�)����5�&QKTѻc3�%�O�(H�.�W���X�Ȣ�2�����׎n�a��s�(��S�>��h��$�W�ȉ��Fk�𣞽S��LC��*C���j���	����:����U/���n2��@�|�ǅ�1,d�PI��P�늋�ME$�����m�}s0a6���5��y���h9����c������S(i#�1Bcr^�C�O����&o�4Z� r�[�������T��:�[m��7��� �iQ�Q5����8C5>�mFJ]���d�0�|��X��`g��z���Ŧ&��B\��xϳ�&�~v0+�����+�^ǸD����XX��j\�կ����xI�N&�g��l�����70X��jG}<��#�>�ruQ�)�>����#�IT�.~u���"�Yĺ�pcy342��j̬��e :��*C��w�\�j���xq��"R�@&SQtuu��F4*�?gn��W5a�����1'l6���vϯ��j��L����Z��t�����-J�RS��PO
�0�,�G��8�pu��y��e��ieE�E����GK��타�m"G�����c��^��U�	����[�q�B��CN����kh�j��q�(�����h��5ۛ��]��?�Ӣ�q�gQ�f�9*�S~�P�BC>nM����y��[�6�h��a�}������l쑛p�k
kE��=���=1�"V�gpmb�²|ߜ@O9(��r�}vtv�ʕ+���=<�H��Y�e���Z��*_�K9�-^B_&���UZ�9�{˗3ri5$���\�'��2�Y�U��{V�����V	Y&�4ED5M"*�Sd1�3���(S/Vu{T��b��9�(k��aՊZ0��"�~��LZ��|�.1����o�5j��xK���5c&-���8DYu���(���H#���:KqVB�Fr�����o�k���&D3�-���#T��5�#��Ҟ
�T�h?h��?4�JN�>N�{�G�nz2KG�n���������~>�rZ������S��U��@ΰa{mfK���������Zs�v%����od4�j8QK,�"K��;������J�t\�d�dG
��N�|�(��24@իi�J��]����~� �l\�P�W�a4+7���Xp�4�f��55z�3*Z�$����ݩ�nF�;�Ӿ�ʾd�˃�LH�M��TD>@yߐ�����#,jP%xHq�ʦi�}�6<}��طf=��B��n�L*��������}��}��;�����Ȩ]Ww:�阭�\ ��ȹ7�Xk�+;fnj�b�d�LV�Vp�[��6����'齝�a|��YV�g���,���IH�9f����O��#�l}�ܪD=N۳j�>�L��\C(�
צ2m�.�7����0�9�����V��<�V$E[n'8�+���{����_,��s?߰|u}#rl�o��Z���/�V/�k��ʍ�:MC֨��Suu5:�n���
nq�$1�K&;�I���E<A͠Ϭ��fJ'���͢3D,���GUl!&�������!�-F�  E�IDATa">�Qlj�_Yu���ڃ�k�bfF�t'$�
.Lb�ME��Z+!�Ok�z���+���:�����!�<b�2��A��7b�gE���(O!%Q��y:��5��H�/O�).��g�a�����3�yK7n��|D|	ܘ]@����� ��w�3�jAf�g��qx}=��?�'ur<ys��Ө��H�]��ׯ\C,���\@׉��kt�vK`��>��]����U�Tݱ`EnC"jA�B-��rUNPǷ����(�/.Q���45/iH�P[�U��`�<X
jv���A�����=ok�������f�!���ٔ���lc؎]�M#����&�i{Ʒ�Ϭ���"����đ�W�lF;�l�5��?�g4=���s�>#����Ĺ����ӏݛ�b�����Q���&�M�i(�u-���Pu=CCk�u�=�S:�J.�t>C�5Kn�9�q"v��A:
ö�݆��3֥!wJ��mKr�sˋګ�r�������I=\�g��ؙ����?��/~�E��7p�ү2���&��#�.ެv(�R}X�9����ϖѹ��.�`jd
u��M놱g�.�?p�]�(����f�����L<QX�G���s�l^�kzP%��Jw��0�X�*��ƍ�	`vF�Vu��M�,�~��L�QR#ʨ&F�y�Ft�gZ.�X�*��������aי�C�Kch7���Ps�����d
���� jt,�ۅ�"e���?U����9��i���
lE�@�A��	����U�ʳ�[���0�_���9�w�q�j���Z�-OQE�4�v^�uI��b&��ۿw�[픀�`z�ĵ���ؼ�9
�tR�(<q�K�ҹ,Ϋ���.��2�	���q>/?��$�p��[���U�cz�f峇]��)$bt���XX8���2F��I�u�U���j�L�OOO6=�6��2�4Ξ=���n�ܹK�-Yz�5WӀ�d���#����u	n�W�p��n�m�N�ߺ��;��ѩ���C����^É_�;��@g�L-JD���'_�c`�������xf�$7M:1L\C��`�[.;��+)��#yeƍj^�=�T�F��I>X�T�V�g��M����Uo��U��BE��y�]��#m�琗�2$��$A�c�rU�ZU�LC����ѦX���m��7x�\rm��mS[uV$'	5��m�N�
�/����o�sZ��Q�����6�	�1��-�Iq�����7%~Ɓ��J+3�lT���$e�I^�/r�|�o�vot�ќ���u������V�֊��ۍu*�T��ʐ���[��-,9-������dÑ3���7ߞm���[���4�s�)|�[+}��k'-<���joS33Zw8�[m��V�C�U��Ӻs4��,.�bR�����>L}�%�pӗ��������A�"����Y,��X�Y�t��d��K�������Y|~�(f�&u-���o�>��u ��N�H�rl;t�B��K#��!TR1�U$O�C��/ҕ�3�*�o	�SW�}5z_]����T$j�Ψ���%����B<�K�s��tF��`���Oo��b�C�&Lg�&h�֊v�]��bfF�@z�Y:A�M�zj��R��!ZG�
4k@3�5	�h�H̮��L�C��Z��
6Ty��A��V(Ati�:Z8�Y��K��ھ�*V(�E��^���;&'��Ͳ�u�4l�\F�l5#A��<U	�����Lkr���Zx�T���*ʄ�B�� j��uI�01q�J������[��f�gTY�`!���Vt�A]gZ����8/KrA��۩�Q��U7��C��0^�_9�c# ��Kx�2��nFT���|Md�M������73C�ɍ���`�*�)��Y�����0�ۏ�D�y�j��>}�:��SQ�Y����O,�2���ze��ߘŊ�S��v�b�V����e\Z����4���/H���(\������W��Uרa�&��uh�%�3��)�T�ȍ�+'ͽ�3�Yb�4Vˢq�S	z�21eل[m���������QD��q�)�Y={n�kZ�Bs��Tީo ��xs!#�f�ZR|�I񬃪[�N�Fl'�h5�{�J�Ҩ��/�,��+lUlT�s��n���jl�,�R���~�QƊFg�0Y���B��0ZR÷� հ�55ܺ����+:�+�U�:H�����r����&[��޶���P&zd+��ċc�eA_�&� �&މԠ�A�2��f%/���oז7߽Y�2z��X�*K�N��Çn(��w�M�ܶs�ޱ'�8��7��Z#�]H 뀓H"�ߋZWWӳXM㳑��ā��Fέؕ��<y!N�:�f��G>AGg��\1�J_Ό���Ku]�K"u��5���X-�����=�&��<��i�&�]ԩ%� ����YI�t6�.�Ȓ�\�3��BL�9�&��2�T=�iN�n�u ���wv���ZC�ng���毦�����:h�ZU� :�rPb;�������Һ�4�h���=
�f�L�ʧs%�噐B�ӑ@A�}�F1+������k8@����*�P�"
W�kA�Q5Ӄ��q��Jf�@��H��ѻnǞh�D�㷙�o{�6��-dXT��h������$ח<�Z��R�+0_O�EՍ#�Z���w�� ����#d�`�Oo=�(տ����B(Q���� ����£O?����y��Kt�hG����rS��w���H�qz~3˒�g����$ZWj�n,	
r]��)9 K3s��eV�kJˇ�ws^�A ~����L#�7v�J�Ea�(Svn�+�5�̓�m�C���Ȏ�X+Ф,�P6
b�-��{q����+���Ew�ˋK��U_�m] �cFu��"��A#U��w���SE�_�0�܎��=��I�`ԷQ��g�iM��~����t��k�H�jk���Wk}Fǔ���To�&`�y�r����y�x�k$P�un�^3�4iϵ{�9����A�b�gΆrp;۠Nh)		'��"S����~;hV����K u��E)-���N���*�M�Ж�%_'�*0��&�Z��c!5���u~���ގ��~�"��\���K�f�R�H:�K�^!�t5�ݵ4$cp�%�͡�)�;9�Oy��Z�9�s�8v�,2)��c(ʃ��0�t$�N�B9��<�sN��D�$�N�������z4���oa��+�,rl�h7���~��oуlM=H`�;!Y
���McV% d�4��B�����H��p�x�*��`C't��j�½��r�-%
L��(	��)w3S)9��H�N�F�e_\cĭ��#��}İc�֋7� �u�s��ߓ����s�����=���a�?sVBM}PW�L��~�1��Ey��Rkz��-Nh*��#c�!kus}LIb�>�T76�ۨF�_^�'g�9n�0��4G�*�"7�7�P�Z�V+zUB��a-ݏ��&t�'��#խÖ*H4���1&����8n렵��C�"�.~4���u��|eІ5��,����O0����,����l�o�N�济��F ��
���6bկCl�( W.�襳�+ױ�U��v���-��kp=�۽��noV�ɫ����y�UC��*-H���m�/Xxicc��������j��V^3���q��o
5���@�Ø�if�#8�0�;���6h�y*�Ѱ�F��Q���t39=�9+�<�"��5��� ����>�q���\7�ѱ��>��y�v<�ȣط{7r��� ?r���;8�ɯM��ʋ/�l¿�����/��}�f<t�ضq���R�,�&�+ˣ=~���w�ƥ��Ʒ{�n��p���Q^XD�|�g�}<� bI񤂔#@q����8�9�9N^>�\U`��:��ܷ��������G/^�	+ac�֭x����^tF�X�ݏx"���T����O>�[����2BYh��Uy�'��Mtut�ʕ���?�3Ξ=�L8Q���?�o|�x�*~���[���;B麵#Ǟe�a��Ԃ!{L;i;?�[�zCm�!	�W|�x���xO=s6/7��'��}C-ة�^k�\�n�ȑ��r-nogU��������ZL`[��x�#x��o`kb@<;Ao�?�?�|�5|v�+�ٟ�M�>��#A��ƞM�Ѽ�}՗cl5
[8pxlɱA�=wЪ#=sENs6L>��M���c���o>�Mb|��-�j�C�:9�X���?���e���{�ŋO?��;v#�ۚ�m*#�9S����X�����!<��S��W8�}�.�~����;����i�.�}�}صu�@�4FF��'9�_���ేA<�v�[����5ٌ�2��.RW�1<�}��Cwc� �
�":��صa�߹����b�bQ#_wG
wm݆ڝwa߁}��?�!>=uRh��o����F������1�����{�{���`��zE���?��F�C���]��Vr��|RЂ��N|"iF]b�֮���at�RXsgJ�"
b�c7&t4I��:�m��=~~�8&�Ű%�5L�TC���-�:��
�Y@�F� �9f�������m(џ��Lælk~�/�i�H�=5,d�C5ש5$2�,���붟F�I,��3����q��\��̑V���p9jSg�ҝ���
l�cOj�������F7a3QV����	��'�J�x��ʯ�A�h�e��a�8����?�ә���gK
Aᡎ��bY.0��!�JQ���d�8N������U9�eʏ�^������^�X:����8s�x�\9���dv�`�%����,
�޹}+��+�ó�?�~9,�\�%2�<}���-N���X�e����J�\�4���r�[���^DQ`և'�(�<�݉�x��!{$�f�&��$�;(�+/y�;r����S�/��)����\������M�E3��X����a������`0�O^����k8u����px�3�G�^z�9�ݰ	��~���@e%��bF��@�Z���e�֯��ywm܉����k��>�L�aE����~O"�_=����y����XH���5�a���OJ��2���aɧ����F���2��R�1g�UM��Ŵ����86����X�˯^�'=\�-��X�?γJ�(�*
��UA��B�&I�+��S,�C����AW"���ی@���`�h��%ι+�	�A�Bu13���V�L�%��Q{Ɛ�k���R��k���5�����e�B�JN���a<��v�Ÿ�R���F�Jd,��ݛ����+8:}�^�)���m�6�۴5?��_/���A���Ice�v�o=����'��P�IR��s"yww�n�`�~���ϰ$���%�k��5�J��������#!9a�'~������Z�E��NV��Trj�Ʌ�,�3؜��J�=;v!���01y�/�ED>|G�(t2B��uk104�; �'������?�J��P2�7d9��wl(��3�C˙��6<u�~�+T�]�~i~3����N�w�y�v�
V�kzw`��[ix�bY_���Q��Q�a]w֧����p��u\�t�r/�,	�\ɤ��w�����>��I��ك���U��c^�e��g$b��0�|�i5��;o��i ��!K�1$RU�P��c�����HL����8�흝�-Q�Н�Rz���:F�>�K3�pei
S�<F�+�0oLq��U	N_"���k�t/��zq��je6գr`���MI��t����_^B�m��g�y���Za ^z�[s�TM�(S�6��{���5���n$-�mه��1����ߧ��ņJ�߲���|�j��-�T�ޒgfҢ\�(y��[��taI_ �8��D-� q���i�:~R��.n�^��6�t��U�^��R�\r�c3ѰсYX��Ρ����BBk;��+t��K�@.���]]\8��lه��$>x��H�x�ٗph�<��v��0~�+��y�� 	��r O}u�n߁�{R�[ݾw/J���^%�\z�)
F�L���ܒ}q1NV +�˾81��B����f%ҭ��s����C��'N��Wi~w<�۶�P�I�j�Sq3	@��J�l�C=<4��ˑ��ө���¨?W��Y�åܸnZ"%ryeI�3a�QB��"���W���)")�����j0��vtu�r!���B&"9��b�~Z�ы;7��3w܍۷������$�Ć�G�/��&�fq��Y|v��;�q����z���L"��O��T�"e���D�J� ���6Q�%�Ӹ�(/��GUښ,�V�Unof��g��s�Zn] �X�ύK�&T�k=��ms�D<;���� D}O��!���]���VX;-mJ�v��Z6��9����[ۣ�2�f���<n"e��I|�XB�����>0J�v��x�^|�������_nۭ�C�B0�Ԓ���
?=�9����]#��б����<�ҋ*E@�2�p���ȧ��?�����\���ȿ��G������.~����Ǟ@5��<�X��)zk���SG1�fw�;��^~I�
����M���/���~����H$�sY5}R�ڢ�g�a��ذq��[���݆��L�t��R�K"���}�Ϗ�kĦ��i�a#�$�w�c�����R9�e�F�����1N�/u����B������,�Q���'ܶ	�?�4�~�i,J~G�w��9��"aZ1�槔5��`�%���'9�8֗�{�l݃�P\�G)��Zqӗ���S�}�Fl���?Ae��8�,�qAOS"A!uݙ �D�|9�$7V>�\��%�=�wB���IB-*�2�y�g\v��"]�
����VJy��(:�(�.��߄�b|�=�DѠ��]�Tj%e���V-�4�R�6ӛkԍ,��Y4���7�mJ�}���Ek�d�y��4b�vPV}F�����;d�SpG"@~y�������y���P黰\c2$�"d ����Lcf�L.�N9���0}�V�=2��[��%y���<�����<5.�6�=�%��r$2�߀��/p�p'���w����7���1l�϶-[�'���e���wp��������[�Ce��T�Z+yaw<�û�a��I,�OIp0(�?)�E#8�e�(6�܎�V� �s38s��Q�q������$q�����k�Ѫ'�f$'�*Ω�ڐ��z�A֯��r�����X�݋�U	j��*������>E���r��
U�>��7_Gj�߆��@J`/����Q�uF�.C�l�J	��"H��;񝇟��w(GS)�=�6>�|"��oC	Kȇ�P�>�I��2	��NY��&�1C�䰯���,�ʬ��s����,a��H�Nc|�����C��o4'ۧ ��7�xN\�oS������p�oš�3Rsڹ@�>՞�"7"��<T3�^I����vGpMƵ����
n"��\D�>��*Uu
5��t���b���y���q��I�wvk��E̀�g�x�>�%���������C������S�_F�l��E���%KĔ�y�ޮn�:ӻ"���ӧ�y�x�~�Cb>��e�d!ɋ�82#�==;����?��)I�4�{�<�/?�<�������V�X{�7�Z�cw�QLH� W�-��op�026�߿�[\�{�aH ������7� ��<��ψ��"'M�mZ��嵧"����Į�a�u���<9!�W"T:+07�woߍ�C됐{�=:7��8�T����8�#�ZX���W������x����fzzq�>tS���8���[J�Φ�!<"0~��&��}j;�Oc.��ؿa7��%T"��hI���a��@�B����ɍ�"��`FZR<�<<6w�n�vc�I���u���<��R5	���d݂#��r��Frog��~�0~��ú��*yE�7InГ��,�*�Y1�M$��P��6�<���6�5�&�Gf�4�l"^���z��r��߀�GdX�L{��\L����0[����'���_��År9,P��T��k_;��6��=��K����g*#��OaÚ�غy3n۶�.^TU75
&9��X���Y��?�=��`�X�S ��GM9����ObϦ����U"��C�4�,Y�3 �ǌ�p����ߴn�ڋa�
��1����J��t�f>6�H�KX�,��؆>�]�� �|6���7�[r�.�~�a<���jvo�>-N� �"oTb])��xU�~�ClX7�����Nɯ��;���'p��U��y]��̣������L\u$G�~�Kׯj����lɋ�.��#�=����������]{j�-��:(�,�a!,%Α���q���bL����q�T+ ԭӣm�P�/1���P��化0��(Z`��0�F�Y��r��-�謊�g#�ֳ����|k���	���U����-��N?0⅛1�����B�V�(Dzt[�4�����5yX���{t�*��ZoSI3���q�T��j�g9c-��ɫ>��4���=1==2�Ub�q��H�P��mވ�z���������CM�BR�bܢ�Il�>V'S��⫏^�'ϟ���4��~C���wq�=�	4�]�8�!W�]KJD�Ź3��?����)՟��_]	,�W�$N�O�� �z�����+�b�ƭrw�����=ay��g�{��x잇�����x6öS��������?ű�_	ԋa�l�窴 �b����t/tBaJdJrN2X�;s�,����:�o�<���ɤqub��� �������s3�����@�o	�۸n3^}i�U!��L�~jn�x�ZH����P�y�=&Z�ץJ�+�M�������=���"X�1�\ �-]�(�l݀;w�Foׂ�unS�&�F���v�z��UlI��^>� �N<-pF��$$ϒ��~��<O :���?��>��]/br#���6�W��[G�v�9����ޜ2L�O�e�6�e�6���qd3�C�.fQ��CHuWv����*4ͳB���xV-5�F�������A��5�\�Q��)ބm����.ua��Q�R��9�f�)�͚A�ܒ����P"����s�3-��
D�B�+��S��p����<��$��ҽ�$�$,�|cgG����r��∮f��ct~VpM�`����ɻ��Fo?x�JC{���82qE����)��1]�"F23�BM"�j��@`A@��N~q�:�����F:����w�)g���4T���w�P0z}��b��nTKt	��p�O�"��á�ø^��5�U�s�C���=�������Y�����������c����d��'�#�KWPXZ���$��"���䉮8�7� ��J�ƴ(4�ۅ��5��:���}c��ؾw&v����TOh�d�CQ������Čc�O8&2��]]�'��3bY���a���z��3uS�olU�� �5���GqW���T�P�n���_��O�^ӠN^WM.'���,��A�QB���lJ������Z3��$�lS��5�U�-����Οy�~�r���Z���|�9&)}'�����8��F�Fr>]�U�)�SWFɵ����/�B��m�R��t�I9?�����oa��lQ��&jb�3�e���
�"�8�%�����;$�q9t9E#��{@!�R?��/�λ�	��@�0��������~�Z���~'�螔�\�W*�1!�݆F��������)Ѹ"Q�|����>�c'��� pO��VLU�#��UC���E|y��b��"�-�{���{�W{��g�
�H�N_�^Qj#X�bQ�!�N�r�����T��<��##��.Ó3�>5uYX@��:��o۪�-�>�L��"!�c�z,�O�!H��+))R�V�m:��m;+mgN�}e����<%Ni)�c����9�U�2�n�Y��}��ag�z4��i�՟kv�:��-�ּ�m�5���QK��(�D�#��qmeR�����{���tg_�2-J٪ Ĩ��{�in�r�*�/�Ӹ 7�����f��#B�(cl���xT�n���F�N܀�8��hg�������r��S���1��p��HHWR�u���?ܠ[�1_��ͺ=]�*��~c_4�R�d\��jd�ɯ��pL��:�;t�s~e�J��$�>ת%П2��t��s�@�2���͆�;vcS�3�7� �A85�u�(�����8vmہ-kע(y���L�߳a]�Iԥ���W�z/N.T���#�FBy� �b"�>A�jQ��,���ۂ�M>�V@J�)��o�pNs�J�jn��nJ�F�Z���\hD!�����8y����ԴFjNq���嵣b�^,����<+�ATÉ����?��+�Z�lN(��X�U�x���&�Ӿv�I�b�	\�6�Apu�ٛ
V����^�'���5��7![o]+D�&}v�+\�Ρ�
c�;��sH�� '�1����)�J�W�������{'�i�2P�6�i;ь��s�x׾%g�>Zh��u�q�����~u
u����~�=����|�"��z/��-E����7QBr���Ssō�6az~�����ѣ���ṧ����o�����v�؎o��<�}����7�nތ����C������?�y�U��!�߻��N�9�yS�(Y-rj����q��w�;�>����r�!%�a�����\��/O����߾�=<p�N}Z�=�����Iy͈3������i�T������V-�U��3�I1҆����9�(?���D	�Z�pa�f��&��~���U� #���F8�D'��H� �g��ɱ�T���+ǥ܊��R��D�N���sB�:4M9���ԟsʃn�cN�c�xBa�Kv��A�u��8��iR.��E�o��v#���e�3��O���H�OZ����<>;�#����*:���Bҏ����{�MAV�2���o�k�fu&�sLS�#(��)T�,P&��-Ć�H�S�NFg���|j�ҿ�U��Kd�I$��0Qs�����<�'}q���;v���s8|��x��/���8$Q��������5����m�w"-�qvn��X*����_�{J���_���"b�{�%|�oj���+���ǻo�����?��g2��ʳ/bIr�sW/�ǟĿ��%��8����I�X�Ј�qv���"����7������0>>��,�3�8;��op�Z	�.��;ￋi����@h��Hؽ��(�1CAc�PqyN�.�g�/�1N*H*�6�s��$-<�N��)�H���[�H���^c�'#џ��:׷��T���0T�J�Ml2���Du	)�D��Ј��s�Q���xC���-
�7�dӦ�׮�^]Qe��_Ur��Un�xDU��R!�b��{�8@
����[k���ŵ�� hZYA�����I�b-��J�G��g>ǘD�F�����=����p߉(4apb� �O"Q^���Ln&I�C�2Ed�0P�nUk�X�m`L���ryɁ��/&�<L�cͯ��f��Mk�m�.L�L��7^7,
9(̧2�<~��7p��%�u�!ܾ�6���j�<\��~����,���,9��C�?<��w���:�&;:��G$z����<��۶�{xf$Ҿ�����o��{��}�<���u�6�����z,LN*�:B�.wO�i.N	Q�έ�S�q���_�U��7�=�4|gf��z��|<6��>� ��R�o>l��ZDRU9�f��S�x���*��:Rd�-�To�F�|����Ji��Y�!��m�z5XT!�W����~E��ج:�V�=������ �T+0�Z	Pyͩ�)��p{7j�V��UŌ�}�K�U�M�,��/ZCs�e]��y���^4
Y����R3�.�06��=P�(�.p�-�7}�GӠvĘW�g�Ґ|I��#�ӟ`L`'�+��9���,��)C�U�g�q�n_.Ց`�ܩ��z��yh��^�Ò3���%?r���F݆�?�rxSZ����!arc�j��x�
���l�\�9]a!#F�-�����h���܄��u���{�t:y��?��;��ǿ�~���\X����?��iH��/y���!YW"cA��GǏ�c�ZlߵSW���3qU�nC�p�2V�Y��Mᇿ�1f&F�.����j�櫆�k$����Xϛ��m�vi���w���w��]�p��������������^�G���W�l&�o T7+��8�H��*��d�tZ���7B����fQ�4��Q%�~c�;���d��o	��"�ܝ���P��l��|�pW\χ�"H�h%���Uݐ�U��f(��*$i��D���{fzV#�޾���Rb�޿�=��Wi�%�mA��i�T�0�]B�L
;����$3���:����9�N�A��r���i���VS�k%{���f�ݦ��+9���&������(�_>���.`���B�n�V9�M~!�u�����vWB�oSb,T+֋��"��r9�bnYy�)��h�Y|�J���(ds��d��O�r|GO�2Lr�9�����xfڹ������vc��Lv��O?����'�<z�a���=x��G0?9�s3�wu Mj����@/���w��(�>��cڿ۴�,�0�q��SӘO/aT f|�WWGc��u���%���x�ħX̥���=u�+�I�{�����]YV�7N1��"�$�ge��㝑׿����c�6e�ıc����Pw��Ly,�.H�.����Y�f��8�\T�Ԗ��VA4.8T�}]�=���`a����d����
t�T�g��Zu�Fa?_�?�@y���Gu�Z$��[Ď�Q��-%�j��H�d�8NeT*�+j
�#7�lC�	L��X*���Uܶ�)W��=�j��I��4$0ӛAޛƢ�����DIƵ�e6�4m��P�|����~}U^c�\�[Ы��:*70��,[q̱b�h�{W툑;�&hީa&����"�,L�����kf��� �C>0��8Y�w���mLؑ����i��$�%\���	���<C�e��J�$rX�.�q#�D�h�L�s��p�Ѵ ���IZ��Wt�CV"�&�:�/�w�ʿqY����1*���#O(!�{c�
��; !��؅/06;�������|�GT�|]-�����a�h���ۺ91U.	U�R���1��|�/�đ�u�$�bM����,ў��t���,Q�#�3����5X����!��ٿy+��ψQ�@�'iH&����?�?X���y�|�ۯb���8�ۣy{gȈ9G���X����Jb0�!�gGG�Hꐺ��)�9�ӕ�Q6��v�C(.,d�A�8�	9',�E�tN����Fg�C'f�,7��Pry?�+��V��_!�.�RE�i�c@��*�Zw���vM�d���/b�2����ܳU��W�%f�JN![�d]�!P3"�VM ]�T�:�U&���$N/�`%$?+�q�H���78v��>��6�8�xf'����aFR�!C~@3S�A�]ϸ��
@e+2j��ZS�kbފ��\�E�$rX��b�|,=)ջ��B|�+�����T%,�aF�@'�!f��n&z�Px8�$��a���2ɽ���NEiJu�� �n8F�OE���bItE����e4���Q�R޲��]����g�����)p��%����BY+������S��U}F+��"Gn���uS.zt'S��x�8����ȕ˗�$p���F��aU���]�I�N_��+:�������p��oqqPK����;���^��sW/bfaV�銊��Y���� �%���|KQ]�J�����>�6p�BF�GV]K��r��8�*����`���S#��عS���0%g�H���ub�"����Y��l����h��!ltH�3K���nS�Ny�����0���Xp)�����>�zRi���bC�v1�ne��NX��dK��^g�ً�ʍa�-���"��U��t �.9�ܔ1��+�`Ԋ����ި����<�	�5D��	89�U���n|V�1��7�	�a��Uj6�3lB��{n���tZ��8]��.����E^�T��1��@�f՗<�xD�QԐ���V"=���6�)/���k�%����3���t��n�f�b1l��HH4�I��c�ݏg�~�.����k���ѻv�]���hxQ�]�R�NВ�t��`�����m��^�W�����عu3�\<��y����Y��Hv$�R-���,bV��\M��,Mr�+��h���q�"�s�@��\9�Ks����8�o�'rc�֭_��[6����բ�ƨ���2y�Y�1�F����Ȇ:0�w����:$>aA:�դ]D"�W���zʫ�NKD�(��}!�YAiun�j��)9$&t�;���:��q��UͲo��R�$Tx���#�y>�#��c��� $%���G�z]ӱ��G�%Ս^�E�*�t�^Q��DY?-����s8W�ㄜ�� ǊIyQ=��Ҝ�4�m�g�c������f��"O�ҍ��2h�F���@���I�`ϛ�ڬd�ͨv釙Vj{�@���������)W�"�A�TUV��-"_0�P�ס���  �ZƃZE�5M��I�J!����Tqa�*^x��o��W����9��w`�6���q k�܅W/��~�S%D����`���:Cv}d�F.���F�{�$�;�{���Gq�����m|�_�i���/�I���۰��m���y�n쟸�ү��gOk�(/�}I�1-?-P��z�3c���`��XcM�*�qqa
W�g�����wPO��e<�e^��_HR�'����'�hB��]FF�:O�?b�.k�l#,�X�kl%�(U��s�;�pԠ2�g�U*�'(a!pO�P�#��W�(��XQr=����R	y.E�;Ο2�����M{y!\�m|�a:n9���S�*�}����E�F��]���Nͅ����6)��y�����'����k�0r�NI��v�9��d����������$R^�g�^m�N��G�(6^K�?�6�)8�a���*�^���JQ_#i�+�S�r��}I�֒K$���kK��и�&�|�U⯫��r\�9V�8P8���iqJݮ���@)�w��/���HiI�G��[Ļ��+&$��{��c��ѳn:�0!�-+�M����g?GlM�����qijNo	:;9���]m��⪗����u�ߴ�l����l�<��utkQ���s��C�Li����.��iq*.� !A�t���q�A�y����Al�����?)���&�X�
cZb����q����P�<����ɹ+�C��0r��Lut�޽v�=+Dl$5���5a6���)��c���AB��t�I6�f
�t�og�7WZ!�o "h�<�m_�6�PM�I�nԬo�'�k�Vq�8��V��̊[�<wYB��9tt�U*V��Z�g�1QL#e%=�+�Î]�������V�ޏ�o.�Ґf��i���:m�|9������5�fߥ��a���5B��®�X�\t�L���(�b]�S������p�VΪ�ȾY��cE��[{�@��i��f�{��Qe�̭�3��+g5�e���6����W'f�x�J]�
Pq"���_�ժQszc���jr`�Nو��'u(�ˋW=?Մ��0�\��]���!�D��1�}�?�ed�<��ع{���Tn_Kze	o��Μ?��3�FA#��7�{w#bԣ��RS
�BǍ�[�R���m�?�1$s��
|��[��
͵\0�b���*����:t��ZB����:l�s��u4~;�g9��[�`��1BZN��*Ϙ�W�~YR��>�	�$+rĨf�R�^�M���Ā
7h#e��.��[�|mX���׶�زK��}͛a�[��#���`70|���\՛�|4��|�U�����JH�is�h�7��������׾�E%&�f\�H���A���'�@�ٱf�֐o�0��\���o�ip�B�:�A�S��dʭ��)�����5L�{2fF�X~`K��E����5�z�Us6���;WKS6�}.2>ʥ�ڦ�����0��qL.�#2�2��^�DK�%,ID�{�sP�޷�թ�m�4]�53�l��׷�s�l�u�H�c�D��ZaP`�vD�	��E���[�V~��ۚ�T44%GϺ��:��*� ,����͵��B��=4y�,���~�雺8J�ϐ"�5MO(mAH�z�i��l�u#�a�=�$�~D�A��3�`��m���Nٜfu38�������,�7��>V�d�Yx����?�$Pv+6Gc�d��9D�;�і[�7�.Z��=�@S<��"�U��Y�z,�k������lBՏNIF-(�ߓ�C�/�����Ltv�]z�T`�Z����[rU�̞��';���zM�#p�ة�L��tt&t~R��kIx��@�Ʊ�p�/�^G5T<[����k�"�o4�
͙�%��ɿt���m
d<	��:::��h9D�W�Ķ,�ߠ�U��5V�#���V�D�����H����ـ`�]͡���:����*o�0�Ӆ��Wb����]b�J펊<E$wܺ�F�乇T����*A2���S�}8J�+4(�ĝu��CU�L��v�o�|���ө�2�Z��:��rx�J�-f��3�&��뺖�6bJi�E�i���Ⱦ@�=A{���BE,�|������#SR$E�I$�x�]�-�ʖtZ6H_�y���Y���{�P�5NV�B�l�?�+���/Lє#Ӎ ,�p�I�C{�O�G���':$Pf�����S�1Qo��t���]ŉ�~�P��`����R��)�RaR8��O����FgW�WI ����&3S�9�N@`�S�襞,Xu#p���x�}c��n�(`�|��]k�wڙ�;_���@M��z��lk�Ŝ�	��A0
�sM���l ��E�S�+��I��x:���[�v)y��ã=����k�^�/F��Ν�x���P�W +=@�Q#cM�NO���y:���N��lb�d@E}�e�	��@�A��I�Q��^�:���[���0A:G�{�T+�M�Q���[tw3!���ġ�8�|H�l�{Fa��M�(]�aR�OQ��}���>�3�LE[����ʅ��ˬ�,ܿ�rD�3�>0���=������%øں;���@������-��\�<X���.�ן����c������*�_���-i\k#T[ ȴ����Q:R��'�+�=zB�5�_GϮ�������~}�i/��`�!D�u�>�d!�������jǡ	�|�wA,e��)-7;`�5���4 �|�"Ԥh�,*�/��^����̥�_P1�~�Yڐ�	Q �C����,Q�\�7n�l�>�
HQ���6љ�siiQ�-)\9���,�1U�gh���g��ʆ����[z5<ƾ�+���w^�V�t�u����F#�i{lC�W��[�s�ʈ�n����kD��I�Z�Ќc    IEND�B`�PK
     T\�,9__�  _�  /   images/05c4396c-27e7-4cac-a4cc-0e5db7270844.png�PNG

   IHDR   d   �   _z�=   gAMA  ���a   	pHYs  �  ��o�d  �IDATx�t��e�U&���r�����s��,�%+Y���0�l��Y`�]v�g3�.c���0��o�Y��5Nؖ-Y2ʲ��V��9WwW��z9�w�~���}�2l��z�������?7������éc�7�U4jM��`Y!x��
E�"7�aX�0��²=����<����.lX�����mp]�W��j1�ᆅP���]4<<��9-~����9�s��˞�s��M~�v��bv�okO�iK�i4�����<�"�����h6��ü9��G����ؖe����B���]���*	c��\�7DBa4k<��k���}�<��4�5�s�9]�����͆�+?��^��&��U���E�r�f�+�P+xK Gu��POW8��������<��;�H/̋��:�ql���aty6��%<�r�9x�$�U
�B[3�F��q W'c������F,F�J�M*HS���Y�!B�r�r%��e�\������N��M�9��z�b���m*�H�h�&ޣ��P�����a���"6�m�Dǎn������J'/����sq��0lYQP�Ҕ���G4��:��X�dx��R;�(bU�&�iK��xx �d
��2��֭.p�
��Q�5�r��fCԐ�2�2�?����A'��%�Q�����_O<��]�DiށS���h,R��4Fu<�	!қAO{�9ԫeک��JLAq��'FMLr��2�92�ƥkX�t�k����]��R��!�V����79q4��C��5�����9��!>���Gp��{W�R���'�o�u��m��X���R9��;*jQ�h�ۑ�f�p���8��:�R�Z�Bǖ�0����t��ȏ��r~�J\]�JT܄c�����y1�(>4r;��}��phP�&�xOǽHcm�����U^P��ސh��k�hg$E2�D&މ��˼�&�ED"FI��S!��c\T
�'���u��UN��:DY�E����#B7�Vb� ,��&-Ϧ���s��D �dR��q�tw��$Z�Kk\���7ӿ7��M�;��ཨKo��
\�g�Y����<�7���T)�^�^�U�R�'��lĖ�?�� ��~jM�B2���~���T���y=�k��'w��C�p\W�]n����L�P�A|l�Q���L�I�
˅�.��^�?L���*ں(��yT�D�:��.��
jI�<�"\`��	�c\�T(�X4���cT�NK�o�I"LY O��3.��@$l�y�MG݈hqXR-�a���r�\��r�B<_�
Ӥ2!�@8M�Exƴ�b�~Yt�!q�vȸy�@��n�� n��P�u9�'���7%��n�Îe|�ZQ�g��wv�����,b^DM�I_!�roG'�wS�j�	�����W����\�
4�.�֋�7{~$�B[w'�Q����jCO[
�|WI+�������<Be��1��u
v����G"~�@+g�%����h_�p�>l�E�q�Z�C�$�5l������(_�@�R1d9�HmY������X�Y�4]Uv��$0�َܵ}�*���q�K��.��(]�'2��B,�����
�ch[���ҧ��K��^p��F5���y�0O��4�a"���-j��2X�Rmt��R�N��qT@bʑH�h+�Ʉ2q��tcyau�o�����(��!rykg&�lQY`���d[��"Y@^��8=�,���+_�P�E-2V$,B��Q{]����9����^��'��}���\U���C-�2>��+����7c|b��������H��#�[}���bˆ~l\����U6�#�PSc���+G��ὓ����Ξ�S.��8��F�V�R
�UP�i*�+E��þ�]&�y��5jR������嗢fE�(�ՌcԺx2������<�R���NLOM�\���ʕ9TN\�U��Z�4�m���
E~�{���\\O��V�,�F~�a��A���W%^X��7�5(C~��ˢ��8n�i�#VtX�KS����H����z�m���4���)��4��Vp���9�7x�z�2L�����d ��4�S�Gi%�N3� $�͖먊��h������O^������~�;���涝�'37F�f��O��T34������;ۻ��сř%�P��d2,N͠I�KR8�\�ӌ��Z@ط��MnUPO��PkSdcK<�p!!Ͳ�`���f�kg�PAY����
U��X�D8�����yĊb�Be�Υ
���rxM^;�w=t7V�Q�WU�|���׮`_�~t2��~y�٬�i>�"��kgq��Ѯ;�W�F�p�@S?���R ��\��h��%�\��>���{������Bh�W�ֵ7���^���<S3�D[52�_"E[{�wuj~{g�mI,MN�����-4���4��m*'�t!$�'�Fb	��H񘾯J���!��!1��⸊��Jdq��(���i�#�'��bؑ�
W��멅���F)Ǝ��/!�\D��46�ވ��I��Fz������0������ƾ�a��Ha�k$��Y�)>3U��Y8��u�.����T+��vf�H�:�y����@;���>r�:�魷���EB��$P.-���5\���;����j���X	�϶jm�P�[���$�Y~�dD�!����vd�E J��s�T��* N��r���)Dy_�?����+$1����F�T(��X���$b �hi�.^_`�r�j�XJH`u��~D+!�E�B��hE{���RX��"�4z�!��#�v=E�a
D���AO�]⃂b[�d����n�J_X�E-��P��7	%�Р?�f�4�+k�2���o��M��.�6� ��v�3�R#�,����� ��(Ht4Rפ��DOn��z*Wc��i
Pb���0�V�y
�,��"�)~Fc\��k�����_ p�v��baz]�(NOW��k�%�u����>ѐ�Y�����,�U�HT�J��x}�+1䫍�˒s�mA"�e!�_���pC�.b+�e��TWW��9�2�4����6xe�4U����0.�z���MN#$��=��/a�J�io'�$�`L��/I�d�����5L�K������6�/D(Dҏ�J�Ҽ����=8��KHŚH1Ve6o݁��T�"kY�,ΡT����m*���ID����V*���Pm8�;�|e0�-�LИ�6����au�0,?53[��?��	�s&>I���Hj�(��"��.�{w��W�R���"���
���u|�.eŦ�[�:�M��6��r管A����]�|_c��Uj���I�o>������y�8�M�nx�~��&,��4��A�ؔ�A��2�5á��F,ߊ�L��bL����^:��ۋ>������46�ڏ���o���G�V���O�m��<�Hк,�*�(�|���]7!�ރcog���BK�Q�".г�]5�)��Lޭi2b�Q�^������uO#���$j�kWtAm9�E�ݭ�0�Obh�=�D�����v��s9L3�������_�<���O�X�����Yj�E��i��?j�����?��U�4k�/����s���E�^=����%I�0���oGi��#o����V���U��&����'�\�/���/�����[���
F��׋vX;1q�+[.�і
1����>�n�n��(k��1օC��E�YqcAVA�"Uc͆�[*Ek��oI�)y?M䫑�w ����^aW��7�od'z�}˝�E�k��Q�?���0@�T���7��$��;��ŉ�ݴi#��nBs�7EA�{��p]Ywo݊�|�޽�@���x߶��M"]�˲�m$�$C�������a,PcM6��B�OF-`�$�<��O,E&𳯷C���JK#;�&�E�ԉ�Y����ҒBR0�+�Z�$�_⸓����j+EnMY4~�Ad����/(��9w�4����� A�Mz�D0�.j}�aO0��@"������ϸ������]ѓI���m���J�A�H�X����\�8�E�J�(�hEM�%bd�����\�M�H�Vx�ܨC��(�ɥ��&k����ڨ�^�jW�.�a�ܐo/J�L��2�@.�0���
��Z��l3Vd���!�ngPm�����1��t�B�p���a��J8����$2(2�����K�#L%r(` d��S�!�O�]S�К���$��~B��[��y׉�I9K�4S�Z^��Zo`�k�Q�J�i!v�(�X������ڌ�_{�~��!�lvm�XG�=�&�6���'F/����	g{Μ}������1�nߺ۝,f�&p�-�117gj���%9'�Z��m���K���df��P�WTSŅy�/�fL(��t�Uq��Ր��b^���[v`���a�٧5����"����LFG�4H7DY��3U��RȲ�h%i�-�� "�&�'(Q,Գ�5����9Fخ�F�|qr�o k=�<�1�:���f�6�ޚ��$}�#�~P�����Y.���,��5ĉ�k�<�Њv�[��.�:RD6�8���"o�s��hglZ^]U�3�8�B����x_�©�+��#��"v�Q�q��&+sKt�9$B�?(u}sZ&/���z&5{��U��]CB:#�L�/iN}�DN]�,��Zl��3c �����p�t놷�x㊖%v���L�-ש�\�Q��<^!W�ؑ���#�цz��	G�
��ĭy���+ o���
�Y�o�����mm�=�#c��%L�]t�"���B���.��ӧ���.ZĔW�ї^DA��.���v�G�賵LFD"��>��^P\��ǿ�Yy"ӡf^"�q�м8g��>[��bW��l*:�&+�P,�;]ͮbf~��8��J�"tϒ��6]?�Z��`�b���(2�}��{)h=z�Ӌ���<�E�V�V!_M-jV�/�˧/#21�����w&Q,�j]ۏ%�-#��a�DH��_�=>�����A�����U�˖����i��U�H�_`�흼�}#�q��y���~ჿ����7� M`��(;�N*��--���E��Z���L-��N� ���A��`M���ZDg(�ͷ�� �s��Wf�����+W5��M�J�c1����t1u�(X�ku�c�����aI� �kk8v�VVV��u�a\������"~�0�V/���h�)�\�U5�*�BQ����_��-ӆ��5����	��t����u'����X�j�KK�~IٔwyL���X�k��E<^�?),����f���Z�������i��$c��o~�>���`U���k�ݚ�6���#Խ��ËfH&����7��|�q�&-a�#�m�C{��+�L.�����{��}X?��L8�s֑˭��7�Z�5�9s�bɠ�fS!y,qs�C��7����W��2��)h�HbM�P��d<��\�(����Dh3s��Ri�"'�lnQ�R��X���k�BB%���h�C~�6mF/9P���E*�y��c�@J��{���-�Lӆ�y}�.5j�
�7o�T��-��]SX�&N�J7b�-�!j����!tL��2�a�PO?:���_E�L�ߙДu���30̋�2g�d;:�q����5ʋut��_��5���c_��Cٰ�Į���sIM�8��-��Kj5�|�H��z��b6��U.��)0�~W�U\��i�QВ��-�h��c3�9�Cm~Ÿ.Z�V��ڨj��@��-C�`�����ض��?�n;|�:)SH'��m�ѿy;������ӣ��1v�@��VI�M�_ܗf���ղ�-$9X�c��Ht��֪�Mjn
��6��1rA&�$�hvR�٠�kN�V�`I��	@�_"IV�$���3x��F'�jf�!|����ƭ�L�N�h�V��/<�����.����e(@W���7ޠ��p��czf����x\
\H%���~�VM$����Y'�ʆ�I�ϐ���&`G�G(�rS��M��i>�w�|��v�ڍ9^��b$�#������D�W����������a\\Kbv���tϲ��p�M�(ӡ*��ᡝ#8ܝ!ʈbbu?8r/Lױ�_�MpQ�;�_m�e�^&ɨHƷj�=a+$��UB�X@��S���c����(T��]Y�+hxT���~�2�D(�T&�U�-`zzZ!΅_��o'���>�G}�R��m�(���O�#(�� !`-ͦih�,-N]�h�6�iѰjK-ʤ�%�'ۇ�Y\��n���á�|���*��ߏ%�J9���rY
y��݇��/��x����ulڐ��b��g�$pY5�/��/��u�n짿m��I�Ձ=�s8������$g Xi_���-��!�� �f�Ȑ8��2�S��ͣ�܎z$N�ܦ��\.�`V����#��7c�]��� F��&����166Nr��\Q��7��P ��_���h3���T*�e��~�\�ֆ�	���~=]R��S�p�t�_̲5q�5���
���&�����ƍ����[nA��^R})�w��m�a���/QA:��x�K>�����GOc|�⛻g���3��b(Lʆlچ�n#�>����	OB�<�h�i�FyW*.��&k-9/&����g��0�h�b���n���+�t��x�����-�u�عnqU���L�������X�[ jG����˩elݺ�7_�t����TC��<���x��Wp��)�y\��S��ZK@��%�s�}�,��vF�3p�2�tjz,yu��k�V*�e߾���̭,н�c݆a�u׻1vm;w�F_�O��j��7o��/����YCtáX����R!tF��%( ��;9���غ|[�鶦�#�>�p^s����������N�>Ot2��V�`�S!/(���3�I�o��SDo�x���)�.1�W0y�n��ft���R)���I��<Q�������lݴi��!\�x����Zא'�M��h��/'��I,���k�1&�	�9�ǥ/)�H4FM�	̵}a	�T��'�ݱav�خb�Y{G�ZSv5���������5�Z��,u��5�ѧe纺���ײ�<��ȅ�5k�폢�����,��+Y��fH�7O�-a�v�K�N�|erގ�b'N���0���٥��+���c�D3���ό�]��AM���/[h���"�Z$R�ˉ؏Ç�`�N(N$�Z����I]�v�r��&�.���62��B�U:P^}�U<��S�V$+���oSm��ýD�۷o�s���9�gg���H��UA�0�����E��������{��)Ҙi����G)�LWg� 6�O[J�}.�Y ��
/��E�I�=�y��6}��P͎criY�4���t�������oe"�/}�+x���� ����_>wZ���[߭fo^=�?��� υ���Fm5�x"����]Q��1~�q�Rn���Q�{�(�A�>c�J�w����F�a��N�_��W_}UM�����SswRA���g��feQ
�C�7n�^��|��Z�}>���I�ܱs>��b۶�<KK�x��'q����(���y|�{�'�HcϞ��+�҂(��;r����}����c��ۆ����,���i��}��a)�z���'�q�'��#���!3�T�U";�T�9��UƑ��<�:��E��������,:�:zi�GO�Є���2�ja��X�pkdҒ�u%�2��҄��)����M�6cbj
��s}�݊D�t=s�d�ytҊ.��|����'��,=�bD�Ѻ���k !P�Z�j�}rr
���R���1�o���*��h�
6l���K,o��K��3�>��<z���]��c�����B,뼿��q]����|� 鲛�Ը�U4+��T~�
+��W6��W.�b�������kb>G��Z�[�E�d������0J��sgϢk�;q
��Mrׅ7(�����'p�Y����؇
QL���f�h�����ў&I��T��q=���`��Kx�g�#ŋ�0�^�SsӘ�kۺe+�z���c���׏�ܹszSҽ"�F,��O�� ��1i{�1Y0��)Il
����d]���4��	I�xSa���V����������ɓV��$�ȵ���K|��ȪMQ��L��E�~�P�ƕ�$fj��(�N�ǵ�J���'$�4n��\�㫳W��Qtx)j"D��\�.Yy�1�d�si����˨�Vp��Y�g�q�ȫ��w �l��.��0�7���ij��VC:�B�k0�G���(/|mM5���^,�h|V��Z2M'3H�%\����*/_�� ~3�3$�i��j�� b��-Dg�ذ~-�Cۀ��M���3�*�%<�,p�Vk�[&m������J$>H�K��ĢT&��;w��N���ʍ��0��[i-�4�5���.5�Д�*�x�q$�`�Y�2$P�KOsD�:��4���6-#JsͰA6^obY�ܪ��-T�n����n0	1(t�#x������ B�K����O]T7$I�h5�����-?�����˫�R\�§���@��ɓkXa��I�G���&�-�0��SJ���4�.�o�t'�~�d[�.CW18�Nc�|I~I�ֽ�f�^"0Z↴		l�NoM��:H}�!���ƈk��>84�Z/際o�����ɓ'i����у'�z�(�MIiH�k�%wt��I8�Jt{UZ�$SK�Qϴ)Hv@"(�4r1�|1B�Vo�I��[ih_�"���XB$(�J�Z��ĩ�C��t4E����f�vw#G?/{)h�q"���,��6�l�U�H�"�/�'\Z��+Ij�p'�D�TG�1*�L�&�GT!��up�A�M��gg0<<L�?B>@B�6�A�.�n��#JZ�2m��$,q �V��o+�����29�
�����Ȇu������=���k?N�-�%�^k'Lo��6�'IZC]p��"*�RPP���1;�\�ǋ@�Q7�HX��፸��a���<wv㍚V��&�vA��d�C��~u�@�(*̓\Q�V��jTK��<�E����J��OO�붂jw�$S�եV���BM��Q��X�hKb�ݎ|�\e|V]l��122��'���6ğ�g�B����5����EK"�:��tBG�S�2��6�N�z�iqIZa�猩�Hϕt��)ؕ����g�<-D+/0�'��7�T�\e����nڂ����)��?�-�MQ�Z����ş4M�K�݂�D;�iF5/������4����8#uޠh�z���JU/���tY(0�e�۩ )D��
�"$����U�0蟥?��]{�B�B�jB��&1<J�<[)�N���B��ه�شu�έ�*z�1!i�v���\.v���u�L�4��)n뫵aGRB0�9AO��Es]a�EVDe�k���L��̬&5M)	�J$�L٭�@d��gv}y����n��Nlۼ���LD4�o=�0Δ�u�M���Ľ;��\�uɝ���$��e|�d*����v	��Im����t#:h�7g����=Iw��#q�Ԁ��G.���.0���ep�9�^|����F�8��/L�s�| /{�����(�+o4�d���w�F.\BuqŸېL�פIBӐ�z-طh�qBݾ�dX�Y�����Nd6�z7��D�A�i��6�t�i�ҏlv�*Tљ���ɇ>M�]���#G�21����#��������3-�C�DA!�#"7���w�-PE:����z��I�?���Z^�b���-Js1�Y��˖1�)��2�<����2gi���d��M�ƌ���}?>��C�dlx���ys����k����Ф���W�g�Kh$�X�ʸR�"�ׅ�JV�풓
�?(��5g�ݝ��Dm�z������UeJ�Vk�*ލEV�0j�� �:DB��'):�i�]*�>�)���{�y�VEm�.���/��u�ˣ���O~\;E�c��̫�6��5��Aj�!7��>�;�$�Cw���
i�G����l=��. �0_Zc�.�FQpLKew#�Y4���.���)��������M'���6�r�@�L�u�ˋ���M�u�n\;�
�$�8����~<X���4���ݸ������Z����
�oM���_$�w�~BW��h�����\�4յ�!u��4t��H
H��d�\^B���ڈ
wg�����6m@%��S�%��!{�Mt�z��G�p�*^D^J�<�'���æ��g?���	��>���Kx��[H�����M�ø�)�#M��� wU�w�v���;�oKغc;x�+����C�&R9�m��x
E��W������q1�\	�M�ڑ�7���m�;a��k��kP�T��x�*�Db��资`z�5C+�M�Y�1���+������D|�ݚ)�J��V�h������[�Y��ǵZ^쎥q��>��M��c��ps�F��"Z�Ff�&r�UxK�qa��k�tW�vD����@"J����p�]w��s�MF�*֑�*��}�M�o�M�{5,�%���Q~��"����Tt%r_XZ�d_�\Ň?�QlڼI3����]PN{'��$��
�٭X!�OxBIrm2����s�	��:����փ~*��S���mua��]f[A
�* U~;�6^K�iI*�C�U���c�yu�%B�'O�Z,��M���069��Cf�0��=�r:,�i��� K�ww��ӈ�G���ɹ<��6�U�U��֣��HZ3{{p���DNq���	AekYIb���`;ݚ[*���0�n
�k��M\�즍�������ؾc6oݪ�l�I.�\>���]�vX�oۦGF2�e
����J-�+�GURLn�'��0)�թ�%�)���|�"1v�=h����D"��N5/D\Dڣx��Y<��c��}�Eյ���ߧ��;���=-/7�-�Ͷh=W(�����g[�̻��0�%9�Ņ���4��e��������������gP n���VT�����$�%�kd#&ǯ��@�#��Ύ�k���8t3��ځ��|K�
adR��A󞟝��G_�2������Fl�I���3��i��m�����1�������]�>l
X��!��b�h����G�v������f�E�����=ԏw�=���΃�ժ�1y�*	d�V�<���^�SKc��\#��b�t/�����І�HB�-u'.��@����7���c�u�m���&��[�c`>�c�x�՟�D�C_�`A4X`3!l���c/=�h�ĉ���&�O&�������~��S8� ���
d��T)�z~s�X�rx-n������-���Њ~������Ϸ}T�݀����Dr٬Y>�\�pA�*qW�������3?���$��&�W4�\D8�®=.s�����&u�����*<uM�%$L�T��m���$�SN%2��/�6�Y�	O��&��[O����}�W��ލ�'��̙74��z���0�������'�b%��1Uj�kg��6�\I��뇇�G���Ӹ�6�f:FTg!eF�n��?/�2M蒮��ڛ�Z�l-�Pl��+.-�����g-�f;�i��6��⋇���y-O�n�旮�ߒ�����Fb��:�0���Y�\���do(�4Z�%��t2�o?�C�:y�{�nm�m�F{6���C&��83�â\�la���f�tꕪ8�z�\.dF���:�9mԔ���A��������Bx��b.t9�$-e��I����~�Z�5x�*5��Dm�YQi����

D[�%)'�,5�����a�OҸb�m�?0���|"�ʝ��'��!1��vx�6Z���gi����H�ǈ�Jڳ�Q����s��T%*x��G�yvu˗Ob�n�:��=a�Ek�p�nقOG�ѕ�ŇI�֕�Z��W�p��h�v�v�<�����ʼd��@WJ����G�/���s�^�Q�z��Y��h��C_ߨR�c8qZ�}Z'{���6b tXuW�.S��U��r�bş -�*�|�7���K�t�1=Ӥf,���-�t�H�)
�^��
M��0{R���y��x�ʵ���� /	�dv���Y]�^�PW
^&��W����7nį��0R߈u����-���)r��-�ձim���Be9$ ^�3vd;���s��]���2ֈ�=c7[�71�0�P[4���͸��x�"Q�8�ɸq#ND1ܺc�xɆPٲA��л��F>�T+,U?q��D�w+�v�(+����%5ny�PؤH���|=��EI�d�� r������k��׵�͡gv	�=���>�R4���C�X��7�"��Lo��)�]��u�=9��z
��|��cHe�6R��`�ų�M�%�(r�e�S������?=�8�|�ydWJȭ.afvE�));��33���퐆�<-��ދ?~�W0:v�ķ��cp�b���Ϧ�,����O�u*Ԑ�YC.�7-V�7�H1I:^$H����"h��j�Tw&	N�ff��Q���:I4�0����&�ePZ�VG���ͭ`eyU�3�H�ܣl��,p���8�K�HW_�q�*��L�^��ɱ��1�\+�X"���F{��:�Ioѩh�3��d?�4�]FH�$IW�����"|˥���s/`ja

���"�ՍI_���<�˿�aZ���_?��z�p��(�g�`M� :��nO)���.���K+�d\iatWv�H#��������Y�^��ROj@�����4k��k׺�~k��Mq� "�C����k��_��̴n���H*U��>�UR��:���I���'��t�[	{�Y�W�9�������5JE���Y�S�Cj�ʱ�
��Bau
���~�M�����%�ɵ�(��)��~�~n��\��޾>�]Q�t���ŗ�%�Q0��mZGH�R~�܏���#k6�L�� ����5.z�75���B=$�6av���X� ΋N�1
$�l]��"�5#+�{�'�~�:tuu�"��w�	S/1���䡙�����~6 pjR�������^M{�zӥ��Ӣ�T(�P��7�)&e�"W����l���[7��}D���ũ�
@�x�Āe�t(�W
�8,[z_�.������jKX�|/]Yƅ�B��:q�"Y��zA�?B�ٺC�5d�v��
:w�����O�B��72��/����*J�%��e�@�~.US����mp�.�t�$cq8��axET� �ˈ�L/W^ٳt�/�,��իػg�v̛�a�l���G�1�_�� �e�TCʿ��_�r׮���"B���dq���>�X��V#���J��Yްw⹅3��<�^م ����GH�ab_�D/���H~/_Z��N�0���An�5H�q.DD��	�%kk�WT&P�7��v/V�8��S����<{B��w��G�;��g���k��"���"��@G/�.��@odI���n3I�$i�{�l5���o���RZ���r�m��4������L��@�~�9BV�A�TB-�J�W��x�f+3l��I��4W�p�����5܎S}),��tO��!�ߕc6�#��W�=�Gq���Q`li��X��}pzC�����I���?���ߌ��1l��<���������XL�weƖ4;7�G%��/j}��z̭,"�_Խ�N�J�+�O"�sHR�(�]�.SSC�b{m���<�^{G��]�8���q*��5-�yjJ����	�U~��	��yf�������I��m�����^$e�b��d���÷�^z�e�$u~��Ru��ת��Ncv�����f��.��k��&g�3������w�2�rB~�p�n���oǝ;v�޽�Fj�sx�ɧt��4Jh�p�7eʛ͠E,��]���$�������n�\�$�$�"Mm�޽{u#��%d��Q.�A�h�t�K�XZud���sy�-A;�m�z��_�'���	���}K�k��8$ʰm�6|�Oᕗ_!��}�ݣ�[����6"��:}ZS?�R�z���i$Q<�����!���҃,QS�!��_m��Gl�r�8��ɳX[���m�q��Pc���S5c %	�O�*,�,J �LG'v�|�D��]��O2��|�n/�9�l݂��_��������^x�e���+�X`��8�̸U7o�laˇ���L�;x�3�t))�pĐRd�ݖ���f��۠��!cF��i��t ���g}��k������/}Q����d��
��UH�_.�t��Q!��	�?��pwy�e$b5���`y~�P����y5���ͷ�-tVhE5� ]��B�[)��3Ia������|������c_��r��8<�;ɐ��>"7�(i�ЦeE����'P��p��w��x��y�~�:��W�y7��7q��$�񵽈�U,N��=����J2kf��c;R������j1�L�mi�mrЭYVw���o��P�Ծ�(;w	O\%z�6�&w�t����\��ԡ42,FcYB��0��s�)��?�~�a�F�����v�m���;g1�h[��ve��NO��Q�k_�C��m�f�X��l�\��~S�ѰA����Q��n���� �M�mY�sÔ:s,_)l��J�Z�g
Vv��4�q�HH��pR[�&�P�����lmѩ��OA����_ى�4�o=���_�Τ���(�vn��s��k<x5*�*W�06����c~��6��t�A���C�1���ϣM�.������q��'M;%�F�Π�t�,Dԟy%.�m��ߠ�������E������̾A���-5�K~WP#�$�.�_��b�(F8dQR%��j�-��E��O�>eͽ�D͌�5nM\��fftƢ!(�����̃�ٿ���ف�J;}
�M�inS���R�jM	S)b�M������^,S �g�u�y���_©��c��� }��&��*�2疗��Z�5�#DN����h�8[��'S�͛��Ʊj[�g\��lm�$�[����`n�V���ŕa�������uP1ܐ�,q�+�K&���;��t��V"�a��)!���>e�t��!�(��*���ʵ�I	�tt�h�o3z:3X�߃��S�!��Z^�.p��s�з�3��¨�*y��i��G��8��nG�Y�}ｗl� FϏ㩣o�D��k�u!���6����Wȱ�)55o,p�]�w}i��b�4�	�7N���-��#Im�k4��\�è$�6�=<�3��P��L쒔K��%Q�IrQ��jY��7Iz����Jv�J8hg���X�T���+<�b�"IP���<Ɉ�*�&L���2�B���*a�4�d��ct7mi����\��D&���n:�=+�3�6��^wY������R��w���m���|��{�<O�����A�x���E	]�Jt��P�����J"�D��#7Yǿ6(��=ӿl���E&a�\V5n���*�N���?��[>�d� ��
o�a��9"'OI��-3���7a��j5�&힌��Jc�EIhg�t�
����F���KG071���"J��57�:�{�����˞_��4:��T�W���xm)5�q9v��$�"v�ȡg������M������D�jYTc�\C�xM'��� �}�����UI�Ǣq���fDѭ�l�y�u\'�1]\��{�(>�a�r���V�||~_9;��taD�M����P����%������ ��}�u�n,H���	�$��n�۲���Y���i%�^��0�H��P �`d���gU;��d�/4wU�f�f�t}w�ۯ/��q��  +�'x��je�n��	�K�����E ���:��I��ה�,�D�L��)6�F�*������P6�D���2f2yΤ�g��d�_=7�W��-�4o�sQ��ZlקX�;�0�فw�ڃ/���Qɯa��KX����?��cs���>�<��SA&GNǸ������h
���&_ӑ{24M\����X]�rUoJ��@�������Tеh#��ZA'�k��K�dedK\�/����aw6��V���ő#GQe��C���h�c?�������Mɑ��	�v�SYú}@� �e���e���!�"V��3}�hR��O"�!r�f#�@�ә�M�^��I�rs���Y���,��S֦/amqso����M�؇f���^R�4�K��u����:*%��I��?�C<��c&�&]�H*��0�޿��ؓ���(�Y�����ǖ���$������,�y��H���=��!-1DjK���::�J��>lR/���]����m��R��ӺNg���G �=��4������Iwb�FD���E��"M$��Ƞ��#[��a��}�z?K�sgP.ˋ�]��t}�ɫ��3���2�v�9r!+���y�$�KU��$Ӛ9�v}��n+�W!	[Z��i��ݽ���%�d��a��;|���dS��*\Y&A՚�X~`Uro��ԺI��f7� �n:�D�x|�0����c(�3djin�J��u�x�z��edZvĔp�O��!;��T���A�Z�?��,�3I��j��=!".OF��o��L�,�&-�����C�&_m�u1�uu����H���]Vn���:IT�X���c�x3q�\�,r]4SsK��f�q��l6��I����,��j�u��.�`hL��
�&�lm�`]>�a0Z�N���6��rfv}�G���/C��A�"Q�	f�����2!��?t�HM]�	��
[ׇ����'=�<�l���=���\?��%d�����0����C�WV1�3�����:���cXC]�>6������1HwT�c�V�8wN��dZ���)�-�DP�%���"��[���{�y�]�,��c��|CIFZ3w�ܩئz���5��A�z�*(ն*�>��c�(����p�������%���"���g���$?P� m��{d���[o¦1)������g���SI�0M�����t��+GI��"�ׅ�IlJ\·�Ó�:�<����{��������O>��}�c��S��O�#�;w�͘��Pw�N������?|�	|�c�������¥��]޵M-%i�;љN!��Ec�� Y���RG(f����R��ip�	
}���U><<b,�swA>+����$������au�>˗wɜ�/}�K��d��W��U
�����$�xB��I#��f;���wta����sh'6���r��W��`n�b��9�ah��X���m�.'��Aj�]&S�\F<���ƕ�d���L4\T.Na�9���VN^BdjK�΢qu�16���<���ұ�+X9woG^@cl���EBF� ���ꦻ�7��Hi��i���³O=��1�eL�Qx��lh3[X7zJ9uÆ:#��� �_7�V쾡�x��>���c�2�_Z^cd�m��N&�8�Aǂ���`U���Ç0���t��Y߃p2�7J�x��4��Ӂ:�]ʃQ������h�$��M�Ez�1�;�Obk[S�yƄۻ]\őǞ���3l_}�E}��[��T�����J�ԩ��M�}�r�S��C��ɞ
9�ê_/}]eQ��ܺ^�Cx�]w)�����_tQ%��P`�F�`����ֺ�?3A�i�fA�FRo��Lj��@4���n;,G�x��,H�3���"(y��ͷ�ǽ�ކ��Nf�k�XY*c�XEe���Jq:��<l�o�P�h1_.8�
�S��E�cI}��-Ӱ�����R���ė?�����-�zQsM�%̓Τ���@C�zք�X�l�w}�Ѭ�n߃���?��VV��2-/p�ely��Ew��EI�KvUJ���a�pōI 6��w^L�'x>�O ��u���:�CK�f�Y+I�p��@�&;����(�]Ǉ�Fv� ����&��r�eg�C�^&�+�{r�he4zIq,,�I��*�p?��c��	�چ��Y��c|�A�Q�-̯}����/��qa���2�b��u��%�#��d�@��~�pV8����qg�����$���_�|n�<�"l����!��e�E���x�)m��M�e �XfPTOO7100�5na��U)w-�@������E�t�,���w��E&0���K�V"۽k1������8r.\T��.c-�j������Q�ݴq��39�.�'��6���GW�Lo�S�Sښ\����a|�y�׾���:t�����_$ƷӼ�<�mX�_�������.^�ً�I^�2zۂ)��2�ӥ�����u�W[����Y��ds��{?�Q|���qaaJ����p�<͓��;/[���u���`#,y*���5I��4:�V&���c�=~�N����/�PYk>�� �9zC�������gO�C7��;4m.��z�(ȯ$���|I����+���@u[�3��Wi9��v�8~:_Ν��`���'&�F�>�����wm&B����2�ą�"���,U�D�x������%S��M��=J��a�����l��Gx�@�H,��A��ɩ	|��#�&�jR�M}�`;���79.�;���*���B��:ȥQ�2E��^չ�ak����B�7^U'͉e��s=p�|L�_�3ݠX��1� ���b���ݽ�������{�<3*�)O�U��V;������
kE}�Q����wߍ۶���o������Z6�W75�X�����q�?�Y|��R�;�a���	=�QR����z�-�҇^�2�I@![�DT݄����<�t\���i�hq2�G��<����^����Kϣ���B��kHF�N�M��h�sh�R�TeÐkR��tW[YU���0�ܹs��b����彆�)�m!&�e��]���L^N�O���[��<o�
5::��7��.�(s}�M�\�]`X��<�й��۲P����w݁_������됀=�ߣ����$զJ6�W~�(�u�!,QS�׉{X֛���>)a�,M�(� *3E��9K�L�J�#�S6����i�F����$7)�\�����5� BPyEKN�q(�����7B��-,�S}�2(��G�����z�?Ѿ5�Lk�f�Õ�����+9�t|0�ҟ���	��t���y��b�A�H���]����So�L*)�"^i<*��p��5�|������8�uI��]Bq�a���U6��>~7�9&�&�Wp��!�9�Sȗ�'��`+���ğ4#���\IP���g4${�e�X���Ç���d���6u���G���WB�\�D����n��3OP�Ɇ��<���Z�Y��7�`I
���K��K�y��gFj4=�͎T���a0҂��<C�z��*+7NK���?"�	ᮻn�I�cS�x��'M��cJ�F �,ȵz�d�� =x�7s�曱4=����?�����$Z#]{��A��(�7����4�¶nۊ�syLʸ�PI��͉v���
�)����HG��쭛g��~��nA۠_�����mU�$�|��w���5��=��];w�p ����U��!�ݓ9/�Z�z��@�����:�R�%_���dD�j]"��v�"�u�-ڋ �C�+���|����"J����G�-������������P�.�`vqKCVsy��#.���Zrc Ž�k`�[Y^ų�>���
�L��t?���"t��=�ݫ&�]�$7�<�I������3�"!�Z����+!l53X~��FgW��1�-�L��{�h�C9cP�uM&X�Ddܔ�u�V�� d�K�+��o��>
����Yq���{��=<��܌��>�����mM��_�z��C��&�~h)�f6p�?��O�'��.._5V�jF���[�v�
����]rN~�c��������ͧǪW�nIyXL�쵗V��X+�l�4�:3R�z�������2����C(�xf���c2���|[�:��;�P��������B��{[�VƇ����hOg02��/_�W^�[��K}ZKܲc,x�z8����^Ŕ� ��|�*�5MI�\�t��� j����=�?�1�!�'֑0����sod����P���5��dgZS�1
B���,�S�j~I�h�ܫ���##`���v	��|~���Ǹ��h'�g�D��b�Ğ��B�rx۶?��yr�@u���8��c���I½Q`f;�h�G�D��yq�*	u���8{�y�_�ÿ�VeMn��$�H��n�&0�/jB�.�݇?��_������SV����--�D���ڵ�U��ܐdI�5T�0���u��/��y�u�t�BeY��p�z	���Z��s Д-Pc�<���Z5���,��R�=�Z��V/�$̿���L����k޾�8�۳��/�~	Y_q� �`JI� ��-��������ٟ>���q��	�p�©�d˘�����煗�a��A�8q�~������v�oٺ�0���V��U*����_j�O"V%>��_�����1=�ۇ���g{��vl�O��E����<&5��m�f��H��1��l�6nD�$[�$�r��h~@�GIo��$���nӴ 3��0l,��C��j�}���n��0���p��I��C���*��_x���-X�k�6�ɖ D5�	��)�i˴u��>�+���x�Gtvn��\�9?ki)�\�V�����O�6H��z߇ޏ�yS�ĭ����G�K��z���n�����g�_�0��n�[�{ᰙ@�0�`۲�~[�4QXV���a�,g�ܕL��A���R;h������+���C@ ���G?�{�'��(T�Z.ЧZ��1��r�$M0�F�z�f���假�YX���?�khڽ!��3��Z�w��׏��p��<��S�2�qr��8V��KI�Q���p�l�0��jJ����-&.�ԧ��8����k?K����A?����e;�>9����*
�%�&Ii�j��\*Q�����9�3zLG��[o���z$i�2��TXM�Ǵbz�|T �\���1d/f�1����KK�����D�$��T`I�hܟ���Vݠ)O]���E���-�e1�2���,ѡ�����.��hXscf.��p�őhO�u�ӎyi�g*w���X�K��&�h���^aϸ9�y�?�.ܞ���j��p�w�0A��΀i�����O=��agΞ��]�ѿ��k�;�㺎,o�܍A�$H�9J"�`˒,K��Ƕ���Nڑ���3;�{�r���mI�=V����Db&A$���ԍ��oU���w��$����{��Vխ[R�J��ӧ`�qy}W��hL�m��N�q�-�t�9iu�c���}�M�q�:io��[nĻ�����������020���z��=q�V\����ǫ����389�E1�]�d3�&B���4Dy����´S9�*4�K�/��&\�9��&�1�R3�ʼ�^s�W�|�i���S'���K9B�s��ZTsR�^� xP:�/jù��FN���0��0Lm��D��͒��E )����	�ց�@����T_�/w�d�%4g���??	�x�,%����]���^\#��T�!�#�\3,<3�(���H�,�����3j���yQ��7��>�2s�VZ^��	[EH��a0͠E9e��;U���c���Vs.����y���1��5��t�r|���C���=�7kv���V���;C�\���b�"�Vdve��f��QDI�(FI�9�!�� ��M�&34�("J?���1QH�dW��p8@t�<����y�6���5:�v��c�B,)�FQ3:�sk1��dk1��Q�4_H�b�1���GWeJ��@A䂦�q�Y�eX�&��S����)�ZT0Xک���Y�yid)�<�pd\*�o�~s����.��j�6ݭf`��M�[�^h�R<s�(h�ǀ�*���lIF�V��u��H��j�geJBN6z�6��9i� ����͜Y���n�/X8�Rt���q�~�����E���>:��D�mfL�^&%��M�1�Yu�&/�Lph�7#8֖g���i7cm�0%��tXJ?����V�2q�L�HLF'ġ�>x#Ǔ	||�7���K�mَ��k�Q�qH�Y>�Ә�Pb�3g_������E�)�]D����sk��g�'3'�����G_� o���j�����x6�#��^#���\�`t(
gE@�N����}�N��� ˒|�H]�0���4;n^?׷�ݯ^R�;��jpŤ�Z�S>�j��a)�`�z�ŪƻZu@j.L^Cr��r�����kVЛ$Pp��T�j�g>�-�{����O�
���L�����<�}���derAE%k����e�t�y���p}�͇�t3�U�Fdd�?��#;�B�� ��`'��qV\_������n�҃g�?��c�XЃ޾���m��N8�NU,v��tW�6GS�Ðݞ��R)��R��	P�$]a
�p_�2�CX6SE]I�Ģv>�n�Eޓ��W�FL���0�v/ۏ���vlݴI��E��승sw�@��ᬕ%�h�da���"��U7��ԝX\Mb�`uq
�������`f��p��Q�<���7���|�&�h�-
9���cO��E��D��� -Fu ��@5����dx%m� �˰Y��U�7��$CV.)C�v�W�J�E��Eso��H�r[��{�`���Wv�f_�9�������Q-ű
W�����䵯�M�%��OH��M�o���[�q������_�����c�������I.$Aؼ1��N;8��J'�j�4���� lp��G' 8�r���0��Z�R;�'SK���xNs��{6�C|HE0�:����ك5����CHx��T�dnL4�l���u���L��No0,'<H��)&�H�g~�;K��2z����Q�J�ޢ�O�̦f�!���]�q����d*.�����U�:/%B����X�dѢ��|�"/^���|#�a�.]��?�k�։>b6ѠT=��@�>U4��Gn���dw�U��$��i�E�BQ4G�v����^~^�/g�Ƹ룓�ʄڭg�d����1 W���`%hay����Yh"K�OɆ0a.�J�9���yv3f�׫@��W�]5����v%�A&���2ёʙ�:�`��%q)?7��6�=�܃���q���;�t��dLM��-Z<���z��
�������ʌ������F!O6k�&�һe"�Ca\��r���	ϊ����F9���-Ņ���C��u�1�Ѯϡt���/���d>I�vg21�K��C�O��ZB\Lz��b��>�&���T8�U���H�pTQ5��K���rN������M��	\����H<�50��8U�+�>)�6�9g���+W��Gÿ���m�p*����=hn�G��M=.���G�;���0ȴ|����#�H�P����t!�2��b1L��BfN�'���׏�	�|>ܷ'����Z�h�o���}�.���q�u�#�����Y+���W#���� �Ұ� ��$��{F@@�B���
��	�\����e��?O�I9R�=g��,r���/��2"BST�d�}��.i)���Y[3�
��T�X�s�Ҭ�"e ��ԧ�}�Lns��d���C���+*$[m%��z	�d��/_���o'�����	��̊�h։�����jDA&��,��46�^H��UKqÊ���9�mh&�8���"�iHE����X�'�2V�*���� H ��DxrBD4��a��C>�0x��H=��k�$�>��L�p�跘(!�-3��(V�N��T��ah�}@W�T�J�*�sqͦ��L�j�i�k�2��K����J~��;9�!�d�I>4�0�+I�s��6�;["��W���L3�P�N�*��i*��<�	a�u��x�Rā�'1~َH<.��ʹ��:��x��n8B~8qa�p}OJ���.���$��#{^��"L>#��>��+vF�I��DFLD��Y�����'�gɄg�
�JԌ����`'8K��f��$ ׼�a����ܐѯV���M6�z�)�R3}΁�,�.Z���M��1�t�Z�F&S8�~��H;B�ݏ8����3�a����5�����r�i�L%��G����zf���z�g~�
*��МC�akȇ%dǯ�u#]鄓�	�02b�;;-'��h�N~�����d�����
���`\CE���M3)���X֍�H^R5��5GY��F`�d,V�x���@&Z�]jz�Yg3��*�2��0K��	)	���_�T��}�LV^�>��0���ke(�G?�9�X�	�
crz��`��YX}����.tt��W���F�@��LKKULR͚5����,G������v��9�E��mL��e!vܺ�}��3Q����)�5��l�@��	�!��Q5��E&*����v���͚�o���cæR��Ӈ�'N��K<]'�(9�"C������p��r��O�2W�r�o�ćBk�2ڔ��*mT�"9*!���Je�{��8p5��_��Yx�o����]W� LȐ�K��Ō�8��!\�w�^�ڵ�q�D7%*j��!e9�4�0�����)f�N.��K���T�}��?��/��Fz��mގ��-���|q��֐]�Q�����Ub|dLxVn2�V]����'�d�2�����?�f6�Q����㒘��g@_v�ޅC�K��M�Z�I9Kǔ���h���@�����T;�(�j��QR.U�2���w5�cV�c�å�.�f̐I��o������Ɔ��=�t��f�6�(E����S�mE�k��]�]8��k�?Ͷ`�5gpH�N�Y�9a��J<�+��G���cC�M� Mit�_��G���Cpx=�e��WbxlL�c�5u�6د؏���&$5&PKN����[tcu��$�3�&O�<��;%m�z�*,�`�{Ww�R��fJ*��?�Ԧ"L6�ݮzHȔJ�ٓ^v�ja9��(�f�Q5)� ��3Ә'�upu�X��öm���£�|BD��X�7s��6�a͚u��S�B��0��kƹ���YU��)���H�դ6^������K7��מ�'�8�d#�H6�px���ÓHdS�p���vcumF(NI����q�$��4ܠ0G#p*�������$�VB0L=�8w��̞#�e�v޲�˅X��O&�5Y�Ej"���P���x1���aW�ה�(i�k�E�����YaZcU�©��4�!�`�[�J&���$�ϝW<��!9�I�]�AP���6_��vZ��wb�օX�����J��'R'f�y�|������	�T����2��p$=	��l_m1����DiU�$������1I��=�j�.�������ħ�KxQ�$�u�~�I]�_���躕n����/[F�U��a9�����RK��K��� |Bx��M��^l�LTp���LF�]�mܰANC��-�M1�v����W9�2������8m�t<�O�yc?b��r
�(#ndO��e��y���9���� ��nڕP �H*�\)IY��bH��<�R��F���� �Y�^4<mGDe�'	��=�W�o`���T-�b������.��!��v~]搙�=��!RQv�;6	
�%��B���i�=��l:b+��kU�����B�d劕�R!��*�Qű�{v���+�3{�L!j�{p{A�)VEZԙ��<M.�J7�|��:�y���"s�*j+D��B�G��N�UV#F���x���ـ�+�O]�"�y�0��o�LKt�xڳ��b�wh����=��={o؈WżK�̮7�f=ݢ����d����Hm��S�?4!�U'����9�Ya3X6WLЦ������ɦ�;��ts$Aχ9a�u5�?.�qԓ_da�8����ɴ����इ`8���^f�Z�K�;K�]
gu�xq�n8F:��!��P5<�^�)Rv����}(D�t�`' 0��D>�Ui� N�2���d�)B���ܗ���6�V9PQU��۷cq�"l�q�Lf`[̎5*�a-�a������&H1I����J���v�D���4���)��۳L�P��_�C�È<���5LLg���@q�֭��ֶ7mJRg�9tw����L�.r�\�6b�^�㐲)1��N�q�X�c��<�ъ�js��8J�r"�_iر�a��G_"W�C�s�pax@8�UM�sԇ*���}I��*��븫C�`���G�����q-����+�����_��8A�3$q�á"kŋ�
�*���8�c��b��4U�Ϧk�r2�Zn<
����+RQR��Io!3k��G�:q
+	l��^�ծ+X�~�2����ŋd&U������p��\��oc0Jc���ۡ�#���V�\��SC���#�Q�VU#BΓ���}�6��m��|�1�;���ٿb�ꍸ�.�ju⟞�֯ۈ;7nE��+��Νx���q����?g����K
����d�[�ŗ�����w��C:,f��x��$� D�:��k��.}������AҐ
�]+��
D0���[ޮ]���	ZT��J��M9�8�~���f��kהC�}�Ūh$���ٸ��qG�����]�����r����s[Z轓G{{;N�9��}D�/��&/
;;�#(�f	y��2��!��V��%�R��#ƇG�.�����"36��j#�Cz`��1iS���¥���VÛ �:8��D�(��q��."A�r�I8�:�7v��%+�a�ʕ
+�T,
טM���ŷ��m\�xQN�CxDű�Gq��9A2k�ߩ$ԣN�E8�����`꣘MCCyv:���G�2��N;��؃�w[��������d�A��{���g~�>�Y̛;�a���q���XE�#>v�8v�ۏ��@A�x��0p�R�Q2���$T5����D�y��P*8����طkN��>�d�3�8r�0��#�c,:���z�'Z*W�8��x�W �����bE�N��. ��������7m�$��$�˸9�g�?�����v)8q�g�ϛ;_�l�A��I�G\�s����l���;h� 1"#�A8�($���(���:��.n)�PY(�t*�p����,�C��]�"�g�-�I�(��q�?����%���?}�f��Gp�'�°" �%{̈́jBݔ~��������r�T�;֞���U>���,�"�)�c��ȕ�vu�F���/6����g��V$�}h�{�K�̓��[ifY�b��Ξ;K7���O���&��j����I��aI���jJ�O]{Qs�	�^�I��E�S�n�y \�7d�&��!��:fce�J�<�{Ͼ}8{�n��f�Y��Nćx��7h��X���n� @/��Pb�Nd��u6Q���rD�`dMؔwe�L;8I�X>	��#G��~F#�\w�dx�v����X�d�w_Ă�X;�a����n�BB���9����C�\vz���qVN�	ລk�����[o��ޗkcd�~���9�����J�������hJU�T�L���l�hC���y�Z]�'��-S���3��_9!iժּP:�S�1�{���=��s�+�)xm���͘=o��`$G��5����Նe؂,��,�����X�7s�ii<܎�x��-OU[�546\�i=n\�+)����I\��:Z�u2λ�����2k�o��^��d��|#��_,�'co�p��4����p &�5ڗ��@��"PY�͉몮��&�=ｏ)k�8�5M�iQˇ�����y|�U'P�tNC
Kj1�J�9YTV۪`�	��ti��U~O�vdN��r�,���W�[��oٌ�Xq#�S�Q�>;��x��O��Zku
X�{�9����;/����E�����dD��|�}	��T�/.��"�Q
׮���'z;ᵻ�B����cG������A_d� ��l
>gAڵ2�l|d��by�>Bl7��5��"X�h,^�8h����n�)+��R�T^8h�)��y���U��c��8��\b�%����&4��ص���%�֥�����!_q����Ĭ_���W	���'�J�ç�TD��S,�*���99Sr"]�������h��0�ȡzw�Lj���AK����w5:*�碫��8���A�zY+E�����}���2&�9B#�J�ܙ�3�G�߇n���0A�蹄�Ed(�J�v)�m8�Ձ֬��xr�kef�А�Q�2�� �|���i����1����5F	ʗ���y��y�J���y=S�,�g���n����٬FIzO8��$d��jt8�d�5���t�l����bdBKh�q:��nKA-$�a�4��P�f���!���~Ct��s��ac����|~��gXɞFW��VBT�o�	2��a����c�~��+]D��E�i����Bf����9Q$���&t�6뒮qsC'����mjbwO�A�%�nav(�kv���1�)��{fc� ;� sNы`��â(8��dv��2��.��O�)ly�A,>�"x�b��{����nYCȰU�h�҂Uxpԑ�8��[#^c���r���̍g�L^���Gdc ����QQz ��L������l_]5l�I��-i��8*�õ���2�����Y��H3����(8��ӥ�06��re��on�B5��D��C�M١��!��6k�suP��z�)���̒�"�I��OEUu�<��c�8�O/�zֲ�*�dK���_SQ#��O+�iK�,��t��(�ݰ�d�ΌL�)P��Ø;��LkV�&y��s����9Yǡ���j���V���� |j,��69�D�.~H�ˡPL22)�w����9�����Jr�١N��f�p�����kk���B$<������*���v�uMl�;2tuS�*���x*��5�?�v�Hd�I1sV�OV�,j��[+��G�p����Zs_��P(S�h�y�^υ(yq�\R��V�h�H�.�t=�8z�^�|Ŗ�����*-���g6�H!�e�nUd zX}����é�_ID�� Gv�9]��<7�sJbt,�I
��Ў���!V����Mo8�IȨQ��
cB�$�w�2Eܺ|-�����Z;~�C�������R{ac{$_΁\ZUY��4��B��t�uزe��*�� �O�V���Ǵ�8b^�~�o��6���AQ���`v��ܟ�<K�nPݳg��������}d	:/u�ܖ��lV��G'%8d{��82n4�j��i�d���y�,	5�U]�� ������`�ŵx��G��+nE��_.�+��p�(���*^/��/\���y�:��[l�(�R�q���L�\U.��bpc�
�lh�������E�&����=��q�@� $���T9�.I����C��L����𠂨Z�';s��w/�lfb���&��h�M688�.:y��S�-�,"�	�2(��r	��rM!��u�#H�(dH�PKvgɂ����{p�������x��\!p��q-)M!t\d�g��b9�r�]�i���ar�tō>��6�ڈEm��/<�W�}����бΖ�*����y�L_%Z�jQAv��/>��#����K��{��8W�����E�4CQ��d��m�L�V|dŀ-Љ8)�o�_�%���@/F0v׮]��;^;n�+��8�`R��V2m֡��f��zY9S� (�b��cQ��5��#22�(X&�1�����_�M7#E����GF6mX�;>u'~KA��T�M-��*G������?�O��SAB�>=������*��g�Òa��!D�H����uuw����
BN_y�1����7����?>n��6�&`�C��GH�>��� ����DM��%.��1�zd��YI��z���&�Bd6�)���'P���>!��4�h��b�����D�@uU*�~t��N��<�e�Vܻ�nu���ڀ��t\����EZ�?���5U�{�ހ=/x��FgGϣ=މ́E(�c�c�
b�8��)�/:!3(p�y�8z�<J��0M�����Xx�7})�����$�9H'�ࡃ8y�ڏ����Vj��)�|��aBundkx�o? \�CH���x�k�K,�3k☒sҋ h���ȥ+Wω2���F��=�ޠN�rW/���g�?��9b+�)��׺�Y�lb�y��L�����@>�c�q�M;���	����@zE\I_������u�J���5]_2�a_��[��U�UE_�Kg�C-���&E�"pN����M�y�-۱b�*�ٸ���J�U!����ؼi3v�����yU(����X9�LNt+�J]	T���D��0���N?IeC�s*̰�_�˽e���k^3~M�E*�o��`y��+��[P�0��ɤ��s���`a+���7�X� �]E`j^�L�t���ܣ�v�p�م�\�G�]@֙Sf�/ơ�$��D�_?�:��ֿ�"������R]S�&GC�ru��&�f�NaUh�۹��f%TY�/�+�q��s��%'Y���j�kP�d�I˯cR9����ҁ�2ŕ9������5=�V �kϲZtT��&Z3	x&�*�.X�1�mֱlܹ[�K�'E�~t��磭m	jj����q���Lu��+�A�.CZ�H�sd�������UI6���G���h�S:K�V5k�B�.D����\�E�)�T2��Ig6�Q���)BUΐuS�	5s�����u�|A�K�7of65)�D�(X�"��!7BΗ�S|�|X��M~G�j51Τ �"����⹸�e-�3�k���*1M����hG�U4쥼L~��^����=VFm�	I����N`���ص��ټ�Kp��2.�\���5i���\!S�i=L�s��l�0X�ӯ��,W]�N�����`֖,6b0>�������n����]�4�NE �x!�$9r��Mf�������n:G�Que5�U���c��#���Y���
�aeK2쾨x���QZ2�/h!6+2�ت)G�d��m�A��.5S�L�L7oE3�oQ����H���R����(������*��5����m+�3�f��*�8��d�ǫW��;B����	�zfT�:��p�9�\%� gΐ�HO���Ԥ22�8�����c8}�������M����_��NL�������[���~ �+�ٻ��R���;�y�%��}=t ���ޏa�%�����u�8�2d������˲ii�R�<�n:�izw�����&Ʀ�V儩�s�e59�ا�����/��������A̯�`"��.����k7V�X�щ"�QA�,�<��bpl}!�X�eA��=���6��r�o�x11F�*�w�����@��)`[�3�����30��Þ�h���������d4��E[�޲Ez�mKZ�����S�"�]g��m�\��t�����"�^��
��c�S4>A��c�	�/�v91l:�[*���O�a���;�B��,zL��*���U&:��-:�UF]&��>��u�������J�΋w����A�̗f�%s6�X>	��Z&��3#n������U�Za��]Zs��U��h����H���Ї�یm���C��7����~^��r=�#�tv�㺕h�k��"�����T[�yn�����d� �$g��Z@���N9�!���7d�A&tF���S�Iç����S�HjV�j$�ET�(�< R9u%$P�b���,�:*��ͨ��ɵ�4��-�3��m����aX�6�nf���t��(TC��]$­�V��+b4��	Y�Q��%��T-_6�|���J�V"m�b�r�v\��ys0x�����31����3'q��Il��Nr`��� ���z衸�a��.�e,�]n��ҟ��j�����s��N��␅ds��e˴�k���}�ٺ��F �	C�TQݸY�AE����8e�E���>��o�W��#���]���tR�`);�i�h}���E��-�b�0�[&�B
N
��h,B���W
9����̳i�+F]�R���:a�q�u�E�hzr�h p09ҋ�(�z��'���ÒNI����r�4�7���q�.?�ߑ��觃4}D�l,��Z:Y���\J�P���i�&:X��f�_[X�E-K�w��5(�fh�DSxӢ5�DGQ�:�>-V�,8�*��qx�d�K�*�}HF��
��`�b�uqq0���~#�,�s=��#S=����2�Ez�B� �����2�����g������!���l��5[ѶlBs��+hY�5sfᦪ��=��AVj��X����<�bj.!K}7��RY�d6I�L�(��<�
pUd����|s�*m�Ųqhƈ�U+1���(��!�%�^οڥ���d��&S�e`��%������ ˑ8m"",YZ��YM(�Đ4
"5�f�Սd�N]m��då0k�"a^��Cn/J�]d��;B���ٓ�s�>�g%�Q�l�Ȱ���Vc|�0f�5c΂e�ݶW�������Q̪�Ŷ�w ��;��;�xڂ-[�a~m#���HQL�B��,�i�k!Ǫ����i��V����g�������U�b�Yȫ�y��yt���!q��d���n5�=*��P}Ș>\����g��pS&G �'쐙wL�'�N��	p�æ���z�v�Y��_]	7	oؐ���o���P��z~�i{I�NX�)L������5��*Ť�]WOĔ���1<A!V�[;y�D��~;Bu��}�4������F� �EP�lW�Խ2x>�&������v�d��1A��$����Zn)���f?G�ɔچ6-�*�ł4��`����f5IzT�2��7+4��L�-���\ʮ�����29�,ݳ�N*w�N��+��L������:����H�����'��4�)�_�:�"t�n�%[A�#�N���Hz\�E5�["PC�آ�/}xt��V/C�����/��-��~���8��8��{�$>h�i���wc�/��eA��z��+2R��*;��)Cm��.������#�|2������	J���6֝b'����Jd�0�-i*B �b�n_��$���[n�z형�.�%�ߤ���o��Cw,N'�E ����A��+�|$1�h��#�_2�ɘ�F��)�'st:��N��+Ц�������1�v��;ЁWvƼ����	�b/����TD���E�9s��)�[Ԅ�����V�':��b��B�Rzu�Y��3Q��qbqL��&��L9�A���}7ނ5K��Ɛn D	��
B�`��w݅�-��#��o/�K-�|��Λ��+���[�`�����/���Œ���	yKڑ�����x�v�=x�駱r����{	��+���w�8)(���?���#���GE&��������~�xi�;���|����?|��8y��GO�s�~�{'��D�)%#��Z��<�����7-H�k�,��`p<���H+J��v��TA���"�?�O=]E�Ǝ/m�ߺ��!�7`�l}Ỉ��LT�Z�x�*���"����lo%J#Q� ;j���%����o��^��]dh����/QD���=���?~�'h?�B�#�r�-h '���D�� B�
����[�a��w?܅�%�L�ba��LW�t)��k��♟=C0Ղ������݀���bv�<���p��;Qf�?�
d����?���?���Q�@>���<��~�y
(��y�n;|�74��%Ke��dr�OcW�E�y)���.�Cb��56I����f$j(R� �RL=�K	m���
�j|l�{�&��[0S�eAJ$k�j<6���r�D�V.8Y� �d%�������%yX��z@��1��s��TԢ�L�-�7c��5��I�ů~�tt���BǙ����я`��0��ӯ��[�n�}�낰�������8��X:��8WE�g���Q��/��GB�Lg����Gk̙��>xS�U�N��୨���ٻ{v�X��>���噡cq���pϊ���O?����8��P"����?������r����&�N7�Q�����J��T	�X�&{�e�Z,�����T$��̫�*l<��6�~��W�է<�Q쏍Ý���N�5VD��x��_a��6x��6UT�/��h 'ʴnk;v�0N\� HL�,����T����жb9����Hn��_��t����O`�_{�a<��6���8Ȥf�a�����!��V�]��>s!�<�UZB:���$��I��[q�w�Newn؂QBJW隄RD��^������N�/�|EF�Å5sZ��=���n�&&B���z<����:�ӡ�B"#s��mVn�_Yq��̰��A�Z�Q��^�i��D��X���E F�*���&��%����߰�ʅ U�R��3���֬��f�d� ��?u?V̚���O�EP��^x�ei?�#W:���-�n�*E���o��ӱWZ��&F�O�3F�4f�4�/>�-�nă7�-]\.��W/]���|]��Ō��%��αC诛���0���P`׬Z�����>އ�C�8�ӧ��_�c�}��mI:)?x�w�껆]���:%����_����3�K̕�ذc�J,��2�LX��_�í��F���!N�g(�rV+���Q̲����aJ�k�z3����Cbv�ƥ�^��pZ��<��\	�ybT:�6��}�ɏh��=�{?&�����Oc�%��~�3�p����?�ٵ�P`5'��o^~��3�W��?��[�<���������qnƺz0�6૬�^2m���{�*�����<��k���:%���O���������_Ta�I�2��Dw���\>:�#��z�ED�O��6��X��u���v�b�Cu*�)Y�Ђ k�)��st~�̺�j�Q4ó'vbw�ni�G2-VT�s�m��T
�"K�LN�"YNl�ia��L��{m����;w`I�<<��o���h��E��w��{�G��S8�~_}�+x���b�Z�}����/�u�\,^���֯���A���??�#��A��n۾�OI|�KVI������w�8)(-������6j�ǔ�0BGé8b<���L�X�Ek���B��LVr�<����ihJ���C��H�e�r�Y�^h瞉��+?�U��PO�K�����ѿ�l?^?��{SP��ҋ��-�%z�A�y�J��?`�JG
S'k\>�i9xT]<��Z/f̚�����$Ep�����}^��6B|C�(:ǆ���9�>��K�ki"�q���,���C�㩤�N2����߽s�ZQ����SH5�G���uuc�vu��q%�Nvu����7�V����%s�����<�Fp�K~(ΙjCع���+��<w��Q`[SIX�I��L/��D�Ȳ��ꌕ.�t��y��`�Z�[=b](Յ�1E��Pb
� ����v
>�-��Q�K���YZ�SĘM��9��Y�jyq<E:´\�#䔱�Z}-m��]�D��؄�q�;�����q�֭Ȕ
8t�4��3�ml2���s�6���y.�Mm�`�\��G82؏{�S��v��^|�El�qZ��!�7�W�N���
���`r�ݐ��W\����G����<K$��{g�z΁�����0F(��+'�����O�e�Gc�R��i�~���0Rr�CâZ�8�����?g�Cz]P�2l�`�������|�X+�O��|B�|G*�
�w�q3�Y9�]T(� jI��E���"ѩ��	j��\r�;�߂��n�6�`ݚ�pP�%;]$|��щ�Dq��-8|�$֭X+!&�n������n:�d�G2���q��E����w|F��G�1`MI�`�m�t�},%1���J6�u�JzVw��%��%(*��c�̈�DB�%�
(� ��x��K��������(NDN�W��Nd�<ZBK�)�r�ar8DR��@XԸ6��@��dZ/�$������zs����7uOdE Ңy��f�8�F|��V�.KO�$������w0�	��xc��~�ch����	�\�H ��(��ptTڬ/�¨�1MS�����֭k�d�2�{������&/^�|��F])X��h��d�au�d���{� Tb1CãM7}�u�8��.��X��៺�E@�JtZ/:��_���C�y��p�6b�g�;� ��`m^��d%�ɝ�E�y]5S���3�_,�8�;t�3+�ˤ���ܴ�����0ctim
H���~nS�?KQ~�d/�D�bxr.pT8p66 +�4W�c6�}�[�GI����͍��̺�k�^n��OF1y�<������/���őBR�T԰y�}'�lJq��k-6Q���4�UT5��|I�>��m3�1YdN�̹�f�Oe{&�c�pN�N�������Q���0B�$gK�E�j�5YL76�ٱV�G"�����9�"N���L@Y�PKQ�K)�t�ezzc�����,�2GVz�t�NT@��Ǯ�Hp=�!�ʣɈ�c��mB��S+�bP� �Ss����ջnujC^���U��Mbh�p.G(�I]��,E���(i:��7m�c
��Z��PjU�d(&�n��{`�� @l�    IEND�B`�PK
     T\��v�z�  z�  /   images/f814d8c7-8d80-4469-af20-bcf736e1bcac.png�PNG

   IHDR    Z   P8�   �eXIfMM *                  V       ^(       1       f�i       |       @      @   Pixelmator Pro 3.2.3   �      �      Z    `
   	pHYs  	�  	�Ǡ��  niTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/"
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/">
         <exif:PixelYDimension>346</exif:PixelYDimension>
         <exif:PixelXDimension>259</exif:PixelXDimension>
         <xmp:CreatorTool>Pixelmator Pro 3.2.3</xmp:CreatorTool>
         <xmp:MetadataDate>2022-12-26T23:32:11-06:00</xmp:MetadataDate>
         <tiff:XResolution>640000/10000</tiff:XResolution>
         <tiff:ResolutionUnit>2</tiff:ResolutionUnit>
         <tiff:YResolution>640000/10000</tiff:YResolution>
         <tiff:Orientation>1</tiff:Orientation>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�Z��    IDATx��w|յ�3�����z���l�ۀ1� ����$`������I$��FBC(���1��m�-7�K�U��fg����Z��jw%Y�f���>�;3w���{��{����»xW�3y% Q��0���4�z���_�y���d�o:tf)�s�/���y�N���@��j�Y�x�F ��4X�t7  �R��2��R����� >��!�J$$�^h�R�~�<�"<�I��[sw���_�`?t���>L�p�6a`X{W>��:� �����H	�)!��$tk�n$x� /8�~�~�3����:���w,���K���Fd�0Qv ��]l`3��}`2+�����+���*�� �p������ts����')?�����u��qr���M2��s� �d�F��IC�'v�Տ��M����dT
 ���.�i={y�q�DA !�!���}D����L�Q���d�x<w���3�(�����nƤ��k����5i��$��I�/V�#5��Z�YK�1�bj�����C}�uJ���'�~�=�����?�9Y5O�0Я�g!��@�d�;2�͘U�7�͘^{Ǥ�GĔ�M��I�33#i�>î�uS�x�	�J����_t��w�2uN�6�Я��v���:		�Ӝ�Ļ�5�<�y?�'Zل�A�{t��w����Ǆ$!!��6]�a�a�OL�hB�ݥ�%��� O��頾���{���,΂^�FO�MͶ	׫R)PY�;�ze�� ��)I�4�(n�G'I/�p^��3E,��~����|o>�6�
�-���$�e���R=6�֏���$�a�� ��Ͻ�ф�Ͱ��El�� �l���fU�A��OJ]���=��7o���N1a (����u���z���D��֯�I!�r���-	�Ӟ\p��ڋ�,K������һRy�}<���SB
��[�ݙ��2!a`Zy��@QBM����j2Y��@{�]��>�0��:���"��W�$$$��"���p�"���:�������.		���X������θ��n��k@`��%!!1�m�5w]뾘�@u����,��$$$����5�!�X��Գ �&�YӁ�㉧ǺaLa�_}׵ VLj�$$$����w]�bTa`�p��'���A<fZy�A�ZTa�� �8i�����,!�s����������m���Ĵ@�V��{s��"�<w��=a"!!15��G�����<p�4JBBbz���vUJF�@9e�����r@M�ۆ���7)AH�	�o<��7Eb��Z�{�	�N���8eHի=+��1B o���HHHL���?"��~��4IBBb��$y�=:`�0 B�:)����7P8n%0L�<Ι�&IHHL<A���L ˧�5q����V5i�QS�ܒf���I��d�Nj}�D>|Q ڋ�,+�C��s�է�ҕ˫�ry�t7CBH�梻-$ ,�t�[#!!1mA,!�'Ȅc�KHH�F�\ixe��d��"!!1}<Q<�@�gNoS$Fc���?�۔���NZ]��b3HbjCg�,7��;m P"��MJ�#8�,1�p��7�͘��� /<JH������HHHL+F����VHHHL?$�H�@BB Y�0��� I��Lw#$$$���HIy(!!�@Jv		��IHHH ������ �0���  			�A$a !!@��b�rjS}�N���_g�������#8Z��w[G��+1����8q�t�nO{ap��Gk�NZ���ן��%���>�;�M�R�m��� IHHH"				 � ���7����#;;;��:��Ǐ �,Y������ݻw/Z[[c�x� 	�ӊ�7���V�5����N(�322����s˗/��`���>;�f~-�%����y�����͛1�"���m��ݵ#�^{�5 ��/3m[k{�)��<�����-�����Ò�D0�N�>��F�L ��F+��p�o�\����Q�:��  4M�hF&hZ��F+܃Q}e��P�hl���W{RS���Hƀݍ�Vx>\���GvV*�N�m�/��Z����񡱩.7�5�ϳ������3\�S� /~M���F�DaA&��+& P�(��	�eq���@��79
gd��ߎ7Z#ѐe2
3��FQ$f�C�V����#��#Iy��iUhi�B�� @��,0�5h��AO�c���I�٨CGg/���>_0���/�Rm 4����ݑ�b+�ſ/A�1�3$I���mGOg�nyc����%!���1��be~k���a�����'Ԉ4�)��Z(�Ģe0A��BFQ 	���	���8,�_
��� �����2�<,�ϛ	�B X0��L	���ܪb�Պ��cI5��0�� �K� �AiI>� 4�*  ��*
aw1P(ԘWU �jU�3�'Z�����_�Z�����p�C )���P(h,�7n��aт� 4-â����80!���$��~+E 8������h~i��̛	�� ,�?$5��T�~�?�2Z��Aլ�H�9��Tj`w1�(/���5�� Z�vG3��l  ��̅�`D�#��HO3�������A&S ���N�y�����g!�) �)��!��΄SA��â����ٹ!��p����f\�/S���B%I,H���u}$�=.G�k�˧~������'"�g4�<^nwx��xU050!��r�ӏd��,8�a/��RS�u��d��={�<HO3���3�ϔ�����~0!]=�
R  Y�)h��`�0()+��2�a�9��3��$�HAȰ�a�vE�7�R �(���������g�d�@��������w0)�٨�F��V������/5�:5(�
���D��0�@pd�%�up�|#�m`���#��� ��Y��׍t�ͭ]P*hm��.'2ғP[��V�� `�#;+vGz-�³y�u Y�)��u �l@}c ���9٩����}[�.�5����317��,;yIf&���`��Oð��(�� �#0��S .(dpn~cUC��d%�~lk�a�q�Y+�|�|D�������Иux���t��*�7�P��R!A�y�n�� �<�r�xZ���^0E�$	p\���+����N�B��
9�������@�7��À�Q���� %%n�E��9�<�ˋ�l#N/(�E�,�./��R�?�I�i�`n�9�ᯗ (�2���w�A�����$���V��x�`CTJa��A(�H�i4r��zdB�i*�o:����`Y^��,�N������X�(!��N�Do__��eA���^������ 
� �^������n�.L45����k%��k+T�����)�2C�ka��Q�m��!�0 �ڊ �X��� V懐�����;K��\�3�x���hh�@IaXg��h�op�[Sۂ����b�d,:|�	e3�@�ڻ"�ڡ#�(/�I�v���/�%��F+�*g��0L��������*�(.Lb#���0u(.L�r�r[�@���N����`�@Ia*8�C��Fp<�Ӄ��>�H =ڄ���a��fCIa:x��kEpP�66����Tk5u-():�o��V}�A���<�ٕ H==贅g���jV!H�����=����.%��p���l��sf���p�<8V�r@�U�+5 &��I�1#�O�G�f��_݌���O��,wbW�e����X5�g��$�8�����y���1h�ǵA��4>k�Q��yLB�`8s,,z�!��0=��k/:��C%��غ��zz�􋃂�~>��zBm�8���<���E�9t�I��Xm+��
����o��76u�Qd[��֍��nAy{G/�E�غ`9ؕh�9�|��!A�����ۅ��_�8,(������QA�h̩3��51�Z}*
KW��^�%���\^��ձ�[�;�z��~�-�ģ?X��d~�Ӹ����A�YXW �G�X�P](:ZS�<�ˏ�w	��_#�B'�E{ze>��6
ݞ�:��V���~x&)�'M�P�g 4��"3�LF� ��$��b�?^6S��<�4����ȌH�$�sӠT�����w|��٤EFz2�v7ڇ	)�A���8��u�DVRz�9٩p{|hi��I�%rs�������2��
��Z�����np�Q)��ϳ�aBhl�E�
��\8�CS�̠�ANː/�o��B�`�5��H��l��Tc�(�B�����l�} {�~&�r��`�z<����������qтԴ�`�ϟ�1��*����A��14*x�B&�� .+�}J0�����{a�ݿhx�3d脒��G2�۩�=F�������~i�8c@+'V�i~�`!�����;�T��}����q� �i��	T�$�tq|~ d()�D�5��\��� ��$fg�j���X��!�D(�g�����h�L�ax�,�BWw�l/������ )� �Q��^LF-fWa��A�Cj�]���Ԙ[U�G :�#:���Q+1n	�� �j5r������R�E��p2P((�KE{G/�r�XX�+�\���;z �QX��nO2�E��ho�I�X��>?7�� g,
[gb����{��x�P��l]���x��˰}�v�a﷢��ֶ������@Qz?����9��x�C���	�V.�P�����]հ����(z�[����.�  P��ң�*���q���-�@iN*ܾ nx�ԋ�`�A�M���ډ�l��;d����'��xۮ|����Ij~>M�
*�f�:F�+��E��>��������#��?��﮹��7g�0uf'~�"�MB ���K3�.�/��6 �b�滮�A���6��7�g�V����gaw�m�Z�&��`L�ǀ=��U��HJ�������p��]��T#l���4���J��
����	������aXx��AkB+rs�����������R�as������xК�����^w��� 2��%̈́�>OD�a2�@��������X�:%�j%�%\�`$ƃN��^�E���B'�M�7�	!��D�����r��7�i�&t��@��zz)d�'�nWNeee���Gbާ������
[2���a0�m�'1��~A����i�[�-��k���֏�>؃�/�;�������8�� �t�������[����h�?yv�������E�ܿF�9����A���\d2��E=9Z��#������˅���/�)�Fu�c���:�t�5�8k�ZA�;� ����{��g�ow\��|9����@�8�J|� ����R��z�i
�|�~���aA��Z��ޞ1�-���V�Ā�3�j�ry�Qk��3�(2��w�}0��p��� �_p�}HO�����$�$bYx�>��$��#��0!x�(�C�@.�0 	*��Q�e����H2r? �2x}a+̈~S�[ 4��2x<>�F��Z%Gww��6^�lق�b�q����G���+PZZ�s<�����z�J�W��9���{���?G�	᭝�������7^��s�pӣ��%I�Y��6��`8���������v���%��Ϝ�a`T
İ��B��j(i�>Ȥ�5Z��c=fqi.2�z�s�_`pana&
,f\����f��ݸ���bР�݌ >_�m6��=�[;#{����,� ��wG<�j�Z0�8 [W_���ѦA'!=���q��0�8�hż�"�&��eY�;���bÜY�()L˱80hhm����k��j�Gr�Ņ� pB����DJ�{�O�ǑcM�8v7��PR��<ꎷ#b�r�`����" �:":���.������ޡ~k:�o�m]�~#�l'����&��!���������??�g���?Ork � �h���6ož�'��N���������e�0*� �Mz�����z���`��2�Q��6�0P�xX�6��o�>��S�#��r~ĎF���5��nCnߎA�]��;X�CSTm��w�o����|.Ԗ'�rص�VP�q<�FI�y��D�>,n}8Zӂ�5Bw���Z�:E�;-�]hi��'je��u�{���u$�bFA^:|� �k��q������?����}uغ�.��+Et~1}��Z�X��)�p��i�X��;����Q[��M�j#h�+AhP�]�g���-���NC���ܴ��N�jѢE�={�I����q>�����X�MZ�g���J%��s�����z�4����������1��Wdl�h�4��=�2���
73R�(06�z�/$	`��}d���Ô�I�>_������<��r<u�e��k��ۏ���לS��.^�g��Y!�,�ϟ/	�o,�⡇�Yg����)F�����<|� d2YD�3)F-�-fXL�OA�K���L�p�o��㱞3�q���}#�|�6)�:��ɮ^�~Íb/��w�+Mf��A��Bo�������A����[����ގ(����m1�(YYY'��AX�r%����hѢ� ��s�l
�R�ipY��Ì�$T構���uq�!�(D�����+��R��޽�"37st��~R`�lx {;)��;Ҍ��@���=�'����?�w�n�jÆ�&�����j9%tp�g����<����/������*�dh���,~N��&##%%%	=���VӃ��T���o�?�C�[��?B���i)���h���7�ũj�^5#�?��7x�=�M�L��Z��JSBUb��=V�����&e�P�R0(d����J +W=q+��v�@��1~w����[�M3+^��w��H��/�����_>���d�P(���iʼy���\sk�E���Q�!nb�uz�vG~�^�[qF%O-�fo؛P�,E�O�;	q���+�h�PD�
��<��19<L|�4x��k���"+��s񷍗�o}�Mם�m�#ŋM���#�XC�|���>$N_(��B!����ۗ��Ɋ��B�N�4�)|�"����M�x��B�aԩ�����4�1		��9>�Q��,��Gn�	���iԴ���k_Tc�o~��o� [��a��ތ:`��֋��߾K����qG1�8=(+����Z;����t�E�\=�|t�8Z&)� �SOà�>Hd����t��1�����#pEW4#w���jhTw%vJl�iÎ���~�����I	�&!1��}���W'�N��qX�;��
��W��!��!9���7����P�O��\��9$���>/�=6
���L���Gc
��AJ�znoI�a	�Xp�>�f�zL3"�����v�����M2�Q87�Ae*�����$��C�]�����4|������ Y�ì䠑�u�>B�7a<��ڕ`B��l�`W�=g�������>b�?�DFm/n������]���OH&p]��㤴Y���`}7^mN�)��`MZ��J�W�܋��Mp"��̀��k���w`�r0(%�� ��%b�:N��Gz�z�1���nl��̬�����N�
T���@F�fڵr�x�@6�;���jvx
"{�^ބ�;p_
�ӈ�7��7^j�C��o��i�"?넹��`��T�&���,8��HX]�C�׺ǯB�$��vcݦg'\O;������� p�_xRj�7���Y��@B��b����t�?���hu�ǟ>�!2���\�	^n]IF1GN��$qz����}�G%?�V��է��n�B>r���O�e�,�uH�D��T$�L�<T��sg�<T�eB&9u�N6�E�EчJ�+�
���1�l;>i����(ָp�ܤih� "Q�    IDATĩ�\.�-�x�`�Rh.,��d)H��-����F���`�a�Z<9�-t
��,f&q0�8�i�� �>���{(��\N&7�a��$��Q���҈����"���1�B��둩P(`�X���
�V�N�V���Gtr������G__�ީw3�ո�L��TQ��h�jY:��v������RY�9�<�2� ��%q��A6�،)����Y��ˀ��0(�t-��kK|�B�&*��Nh4P��ZX�"��_��5k� 99y�{^|�E��cG����lFQQ���`6��L�T*�s:���l�?�]�[�Q�cM��4V�%lP Yzs,,\A[e��.3�ɘ����qsU��G5iX�Ϡ4��3���%.������3�[�P�}o��ڃ����@&4�.@R��n=8��Za��$##���Czz��Z���z��z��;�N������6�-?r"�=~��'�k�����"��8;kZEW[�����,�8. (0q�qv0.�`���e3�$q��!:�dU�i?�D����X��8�2?�ǿR�%!7�;��������.���qx0��h���vp�o�la0p��g�d2a�Νq?��GA&;�ddd ##����*�
K�.EAA����^���JTVV"���������㡩����,tV�Ue��<^��|y�?y�=��]�����w
ӓ�x���/}_����J�
 ),�?��_�*yTԚ@�wf'.�0*y\?+���3~~�y��p�L��:q��?b֏Â�~���~��o��~��!/'�TӸ�*1k֬��Z�B!��fTTT`ժU8��sQZZ
�� �ea�Z�DI~���d|�[ߚA0�\��3g��/ƕW^���*(�'�Z�P���ICjJ�B�@��y��ȷ�������Y��ƆK����]�$q��/�-T4��V�C�8\P(����*SY��L ��`[��!�%ڔ���窌J^P���6�$*�2�į^܆d�Oo�O�z)nx�t��x��j���Ƭg:cQ9��>$%�c���7;�(--E{{{\��Z�*�'�y���hooGWW׸��5k ��Ǽ��񠫫����z�p������%>AP*�P�TP��0�0��0��qn�ш�b�ܹصk�f/J�����ߋ��dX�̨>,�o4�T7`�?��]s.�b9n�xh�ē����ڎ@1:��A���M��=��G�k�\Q��+Q�dU:37�� $��0�vV�`U�ܬZ�΋���Ǽ�Ǜ�&��婡���?'/�0ΗG�q݃/�;��K?��?�rB�g�'������_faA*hZ�$E�x<�x<(����㸘�;�$�Վ��7��LEA�P�����|C��j\x�Q���C}}=�����7fpm a=�F�1����Ύ��2�K�,�Z�Ʈ]�b�8��JAW�+�d��0-�i:��/��!�H�<�?	4�cY�P��r��v�k�uƫ���H�W�_?�(�ؙc�FhdepV��kc��G�^���>����
���ּ��Mn ~�ۚ�\��k�zF%��Y����q�ٳ��_ี?���������� �����?�!)�H(V�xزe˸�[�l��N�3^}u����^{툲�:�X���{��������Ʉ��Rp���lٲ�@����/�J%4��,�}���СC��1�n��n���ѣ�(
���(((@^^ޘ����
6����d��00�N�p�����,<����N6�ww�Oo���ל�{�\���(�]}GZ��a�)1s�ۃ]V٧�y���������w�L���0��뉊To��#�����s�{��^�т`8�>��#7"j)A�3���c��[���~���:7��`ĵ��d����Kc�1D���3f�@F�hh�m��N����Gcc#��h"�A��"--4M�III(,,���~���{��99�y,ˢ�����P((**Bii)L&q��xVlb������]�2�umc�醘���Wz��l��gϠn0��o��1>�n��߽���8c��#�w�Q�;���W�S�G{��_��/�۟1��/7*y����S�a�ɨ�c��c��X}�7�T��zV%��Y'�Oz����h��Y'�i��t�`c|��xػ�r�,�X�o˖-��gbE9�Ö-[N� M ��Çq��a��梪�
iii��Ph��Cp<����@���0�����=�������￪i��?}���#�|�B/���H�ޗ3{+<�G��u��@̼�@y9�KX���d��-{j�fԢ(s�U�R�$+eL_����89�Y�9w2��f�� --���}�d{/����~&���cFzR$$z0�bw];x�G�a���k�A��Ğ�B�ѣǦ@8E|44��]�u�ވ����g��:p&࢜�bĿv=R�=����sp���.����#���3>��S�����C��@�Vʏ��5�tuu��ߠ�07\��J�#-.�'��t��b���K ��xk;��g��w/�g�����$Hl,%k8S��wi��$^�P��Z��5J�'�N�I� �D���&e�Y���1b�'Y���\�`��ï}��.?k�,����卾�5��
�J����͸0��ͅF��0��l���k�sN
����\.CJR�LeQ���aP���?�z	>?܄_��C�<�+Ϛ�[�.���,,,��O�}?�la"cI'q~
��f@�犍U�&V�q�$`��>V����Gy
���{n��ݷb�SOE��6��
��fI[>��N��8B��4���*�T
\�ϣb0�bG�#�RE"q�哴�lx���c*ńg0GR�o �)F�e���a���7���uK#���c}$B|�48�EYܥ�ƍ���cw/�d�c��ݟ�������Y]�.�i+�o��"�2�e9�s�O6|̰|���)+�Xѣ�����c�bР(#���sF�A��~���.\<��R�e�y؆Olxx
=��\t"g �	E�'i�X�l�2lۖx*;�b�CM&]v�q���5#�tbMa����'��n��PML��������;� �g��aI�H}M�X��ܙ���n���X��Rɉ�\=�L�!��/Z�VQa��*�Y9,2uB������Ѕ .���.{:��v����^��6^��w_�׾8�sCx��.o<;�p���ǃu�x��D���@_ٰ~�r\	bNuf����޽{�r��P(PVV���<��/�su ������j�����N<� �:����qm�O�1�C7��ay&���+��Ŋ�-�x�2om�a�%ը�E@��K*0rWƪ��h������A96,�/ǃ�6W+�γ �n���x��r,�� ����#�:���ާƬ�h(^�jՉYj�U�:i�,���FZ��������y"W����D0�1�>���6�Պ믿
�F�qL%��n���(srrp��ѓ��)�h� ���h�h�ot��a �ݎ>.{̺�̉;�Ep큛.�7] �׏�����H��
�|P���&d���E��:�I:��=�#�}r�<;�*�Q= �����t����W��<���
�œ�����El��nb!ק� p��1477�ħB����m�<Q����с���eeee8v��)��.�$�qĨ���ۏ����0�_���;���u������A���o��x�L�G��p���w)�����tVx�aCٛ�SG��t�����q;����B��6'%�:���҉^���_s<^
������dQWZ�ۍ��N477���U0h'���R��ҥK�{�n8�N��rTVVFE;#0�Ç���l�̙3�&ƉP�c���'�J2�Ŭ����,�n8 4��0x��ݓ���n
=�����z�p� |�Bc[�L���17�� ����q�*��dfU8ށ�!��j�(��`�L���"8ˬ�r�����<N#>�OG 
�Q6\=�N�P�D0�LX�p!rs�+��h�Z���>����Ç#>��["����:��� --k֬\okk��{�����jEF�H�����W_W�:n.�ſ�����0���yȴ����T�qs���MOL���E��=
�8T��(2�0)���
�{��&�3�Q��c �<$�4�����1~GU,��#����� B!/d���q0tz���d\�G�Ra�(++�'�|�Պ`0��?�|�m:z�(���D�8���޹s'.���F�B�իWc˖-��2qFN��B!7d2�0�. dY�h�k�K����� ��$�����":2�@�ɦ.N�F���U���2>M�p�Z-V�^�ݻw������y|��G���Avvv�騻�	�2���Euu5���F���f\}��hnnFSS���NY?�x3S�(8)���`��C1���2��X�z�����B.\�Z��۷O�>��
�����ݻHM9s�$����eY�߿�����N,�M�7��Y�e��8������_��J������f����9���8��r��� 777jt���
�A�ٳg\�[�bEļ���{/�=?˲���p饗��W �T�ϟ��������hm6���q?��8�a�&�ۣ
���@�"!�(���2�$IbժU�����V+���+�T*��磼��$I"``` ---طo_�SP�<�ܹs���=��F�1���}�g{q:�I��D�����r��$_�RVf2
gd!�����w��ؾ���`�XD�8p ���X�l�`I�H4b�X0w�\<x���:V�Z%:��u�Y��?�9�8�0��/�$X�Z��ڵk�׏m���5���IX0�2����P[��-v(��D+����"��p��KP$�0#��yFn����v�l2�RQS�O$A�hF6j��a�,�d�'��:f��	C�4�̙#z���?G ��u��
QF�4�ϟ���4��袋A�Vc֬Y��.���{��F�ں��,LV�X1� p�\8v�jjjNig���<�#�,�FgW_\юN&*�Ǚ�!�J�>�� ���'�U�G{b��b�2�,�.g����$�\`
by����d�:���=9"�Q�	A1�+++E����n��ի^&ggg㬳��֭[q�%��VTT����	E4Z��t��@�RE�&n֬Y?�!�����~���'9�P(h�����0��϶0#����Q~�4ţ"�EE
��/�c`��Fc
�y�,�,
�LF#Y���x��{:
�½W,��,�evk��m�i�C!N���&�!��*��՜P[� ����x�^<x�]vٸ��YYY���þ}��x����r9���P__w}N���-��h�Dv.**A�Bq�nS(�+!����W_���:�6�
���`�2P	�R��Ǥ���L��y��?�%$X�38;Js1
L6,�o�hu���
��� �TH W��a�8��@P�2����p���6���D�� �V���w·A�����2��T7 -��R�����d���"_ ���CEE���������hooG0��dByy9����VUU��W_Eee%4����������(..�Z��q�***DC��嗧�a����A��u�iftw��ݓ��C1�g�U��k���O��"/�� B+���9A<��\�3�"�Y��!H����_R���Us�p��l��p݊9(�I�o|�]���~q�y�����'��v��=u�F���ǡ��W]u����n��o�=">���EGGf͚%����GSS***b�{,Z[[�s�N,X�@`5hjj�ۇaƌ������R0hnM<�Z�Q�\|�5k�ͱ����h�25���rO�Ɵm��y�����w{�' rE�<Y��>3��'%h�r��2q�/Ӄ^^��ֽu�|�Ux�_���6�iō�惎b�z��T��Sl~�#�|����m��`6�A?x�Ƕmۢꬮ�FFFrrrF��������a�P(��h:�X]]���:���A�T��󡿿?n �^/j�ؿ?�@_7r�Rp�y���|� �]d��H�c��?���0�������9�x@�B��-����
�X�8�&����@�(Ch+d8`[#������V����߹񇋳�'G�l_����F:n��N���ωze�@ЩƎ�S^�1��/��|�0�"8�N����3��ѣG��d2E=M��j�:�.�"p8�:e2Y��N�s̭������
�Ӂ�` A	�c4�՘W%<�7���.��a�s��u+��ŏ��]#��Y���^,|P��G�Y86���Iq�;O>���} ��}��4��
�.ʌCdh�Y�F��*�t� ���#��Y�߷��Jc/^nP���qQ��F�>ށ���q6�@8lzE���uX����θ�SN5b�A^�WԺϏT��Ju5�H����;/��ы/����`B�O62�,@EE������W_Mk�����[aҪp���xg�1|q�9r�b�+MeE�s��m%"���O|�'�n[R`�F�.%I,d$F�!Fi�F(8h�'7��P94��)W��MK� ���KH1h��.įo����s��ˠV�8�ه�|9j^�V����u��i����ɏ�Ѿ�Iϰ-�Xy<���+��d�<��Fm�h4�[��������ٳ��Gǃ���;m��Gxm��(��`0��vw���,�a�_���jZq�Y�F\붻aw���b��"��/�����X��z�GF��)�0j���t^��?�ۣcn���G^�hi~�4oF�#-]X��P��8��1�.��t4v}�&\�x�`�u 8jˇ���>��\����� f��h4����������1}Fo����v$��c��܌@ �����~477#///.�#1a:��1UX,�\�R0��GnJ�P���da}���|��]KШOj���ԗ>4��b�`B�������5��'�j���t;6msv3˙��#�����da	�!

�қ��}�̃Q�I7m�D*�^a}qNZ���-k�@�Q�l�Sߎ�$�Kw..b�������x("�8��Zg�����[R����z��r,\�_~)n&5�5k���f���1�<?�pi@__JJJ�r���g�!))).a00 A7��x�x ���X�p��Gmm��iꃍ��	-v�4✹'�7�h
eƬ��Q�p�2�u��[��}/�L�bn�r����99:><��'�v�S�4�â���������a�I����v��e~��qޜ"e�Q*h|{�l��J�}���X�����>��V|?��'M��3�LP�T���@f��Lyy9��)�v��g�� ���0o�P�=000�|>�v�)I��={����SSS�x���@v��9��]>��5*������W7��g���I��5�T�$��������=��5�v����SE�ʓ����)ٛ���~�����?��;�|�`��G?1�=�.q� ��8oN!.�_��zo�i�&������s��#cF�ME�`���h5���Fz��EF�@8,��}�� ��F]��`{{;�^�h=��}�����C̚5]]]� ��MJJ
��������ݎw�}wB�0C���(K�F~g�:�-A0Ɉ:HQF2���
�zq��"\������x��=0c/��H�UFS<f����+rŲ�_w�K����.ow��ک
Fj�j��آ���e:�.���ˆ�_�q�����4/�fk�ȸ�����L�qu�������A��U73��R��9gN
*�m���ŵ��I�z��xD�̜9�PhB�8�@ _|��,Y"�N��p4<�����ki_SS#x� �\�s�̙���4M����֭Å֡�    IDAT��^:� ����[o�5�	�d=.Mk͇�$8�glDI�H+�^��չ�P"zP�!g��B��P9E���Ǣ�N�Ț<DY
���4����Z?";��wn�8;=��R&\��NF�����)�h�Yz^���6���|Z�T-�s��y`kct�9�|'��ɠ(�]_FQ���d����	"3M��/q�;vLph�$I�}��x뭷��jE�c�0�n݊��tQ7徾����ٳJ�2�K��/D�}��g�i:���C��;��$Ib��(--��ÇQ[[3]�h�F#222������̘'=C�v�ލÇO���3*�1��[�)&tZqOϪ�T�����l�?��M8������UOY�Ud$,��zg�#<z���bD�;H��8�A�����2,�N� ��S3���vڝ�y]�?�>���U3�N]�nV��ƞ��LZ$��X�����={���o6�q�`�֭�3gN��Á?�F�g�y��=�w'����EA�PL��P(!aSS:���J�5�V�ŋcѢE���GWW�N'�^/|>_��r�*�
:��III�g�q��q�޽���JP�(Ȏ�L#YKc�Z,-˃�$ܚ��O̝��
2H��z�⑭���.�V-�b�*rߪ����x�E}?�7��w�L �������0,�"�����رc֬Y#��%r���UUUQ}\.p����f�X�BTx����+���矏���WF�8�رAܤ� III1ߙǡ��	Do�ɍS1Q�^?X�Ý���o���� ��~P��`q����2�r�8�0`9�o�帼4�"����c��YBAN>>؀�>
r�3bEW ��_? �>�활����8p���i�!�]oo/>�P�Y F\S*��������O?��O۷oG__�.]W���v�QWW�cǎMz������/7��y6yP$���mG�=9#F�	!�0 �)֞إ�M���+18x��Ƨ-ѿ�1���|D�]V2�4�ñ�I�SO��w|�#�"��;����7N{��ARRR���x	�B�����׏��f�z�!�`)C��֢��,=�8^|>ZZZ��� ��z҂��!���7D�D3�{0ɫZW��v+�83��!����aE���it���q��^5�
X4f&s0�x��<\Av?��^J4��t�Q+PQ������m�=S�n��u�V�\�RT�7B��l�2fR�x���CMM�$��N�۶mþ}�0s�L̘1#a�`�a����͆��twwm"%�?{���y�}�s�-˶$y�1����!���6�M���4m�~�۾�f7}�4MҤ$�@{0{���6�C�e[��:�|	�:��������Bg[:���=�q���HI����Ĺ����t�0�Xl�X� ���chDK �b�A��L�AGBo�+�͵f�I�����y�����Bf���V��E7�0سgf̘�iӦMJ��^�Ǟ={�yC�����ѣ8z����Y.�C&�A,{j)�V+l6�z=L&�u3���V)����6�"!fL���#��b�h!�:ryc�Q�H( ���n4��@�R\Uc ��'N���s�̙�uh�F]]N�:uM��&
�^v;���J�ᑱ8���I����m~�q���$	,���=w��AEOO>��Ӏ������~��I����l_K�r-10�GA~&F�vH%B�\�� 7�1 �SUM�R��8M͝0�J�R`YvBe�W"w�e˖I���GF��֍�t�6;N�n�֏4�!����@ՙ���~��A"�@��@�T��(��vA����H�v���?f3Q�e��,�Ub�䢱�刕��a��+����R��U���2l7$	��ˑ����h�r�P[[��gφ]�|��R�l��i�]�����F�"KI#Z�B$ F������!
V�C��1H�bp[�Y�'���z�Z�h�ѥ8�X2��8�o��L���X�lYPU%�@���deea۶m��%�c�j���U��~A�e� ��8K���h����E�� * ���N�3ω���Ȏ�6�ʊa��L;��u�ȯ}�� K�.���Fdd$��kƊt#A* ~8݁��A�)��@�sl(O
^�� ���M�J�pS�Ms�e�MIG�_��(��;���_����������!\yނ��7�f;���×����q}ײ�PPP���(��ޜ��{0�R)fϞ}ş�r�����~|qL���Z���L�4��?p/Nz|��St|�<��Ϗ�����ƹ��Bl)��ې��_�, �5�,�<���r�(���fQ,��Y��H\�jE�"���Mxty��u
Ͽ���h/����g׀
�#Ĝ���kp�֟�{�`ƋGD�2����L�Ք��U׆�FC^^��瞞lذmmm�m;v���S�|DFF's����*��qW:*M��/�o�4��?��Po���c����aX���;!����yBl�
����� ,v ��0�eל�+!��� �M#V��m$�zp�� �	�<�^6#����wk��}��ǎx�_�Q���z2 �6�o&�];
|Kbw���|��`,h�T*=��}�v�������O��֭[=�	��dm�^p�M�:G�϶.&'�}�#z�8n�oN�ƴL4�H<��g�p�i���Z����A�rt� ,���DF�gA w�9!���4��\�n�v�t�h�엿zC����z�s�|CT�A=4`&���HX�~P�d��O	������b荾�2`�o�Y�Ó��FQ���1e�H$�$	�Z��O.�C�Pp���&I� ࿫��H߀mUU�g�{��G�V���K"\3�����wP�f�".R�cǶ���M�o�� w�0���,���Ͽ.��o߈�lQ��uQ2;��B����d����9B����Q���]���C�'��_���_���"��T2_���X"�?C2 ���8>xv���`g�ح�����!�"`FL���$��m\�N$�rӎO�/�t)�b� 99f�_|�E�
�+Vp�����v�ƍ���͛ǩ��ƻ�0��jժIQO��]T���h�����F�JpH%E���X)�N���ܭ�3�R���: ���_߇�?���s�F1�MC��&��/�̚�_x����}�<y`v�k���}Ȓxگ���3Ȉf��P���|�����L�����=��o�@z4��Ϳ?�-<��4����<?XV�G��ī]�N|;]���dZ�(h(����nHē�2��̌F#����T*����ш��N�}�7x��}ڞ�e��ft��J̉h��V(�FY�/U}�2�b�@ �r�p};vV5�����KK
�AЏ����U��%T�U-o���>�}����Ƚ㷧(Hǹ~�A����N��pJ�y..�y�������@1!2�8�҃/�7x�Mv�jB��Xsˠ����v����kIL+fdEB�+!��4j[�1jc��$C�:�>�@p���رz�K�.�@ �֭[�|���' ��~��n����hhhmohh@www��|�����t:��� �Ӊ��!�T*�Rm�|
A�$I�e0��*..�	8^�ݗߚ����t�숋"?]͙Z_:C���>nu��?~�t��ٛ������y��Gp��⧷�F�.t3W���3��=}�P��.�u�Y位 �h	����1�p�v���菁sw ^xa�����"_E%	�%l{�~��&�}n�*J3�P�tB!��y�dpWԕ������A`޼yHHH�������% ,˂$I@$ ���0���=��E�eY��q���y���zl޼w�}7bccy�o6��p8 �@�$
gw���ӡV�}x�NgPcv� #Y����ǥjb0h�� EGN���美����x=�ؤҵ�K�����R$�o��8��eB����'��������3Ϩe�����3���3� -ޟ�t�����������}�YYY��ʂ����Daa!X�Ņ�����VEJOO��?� �*5�d2�~��P(x�wPPP��s炦i�߿�'�w���,z{{=.��c�=.Ƨ����z�0�HT)��/� '�?Vs��?|�3^L_f����Q�-\�-���O&G����$�ˈ����P r��EP<h	]���T`��߅���?��O,�'���?�Z��g���/OB�N���./͸}�v���A*����f�YYY����J�� �̙3�7o� �0>���(,,Dtt4��\.��ٳA�$H�ļy����~UB���=� +++�3���Յ���+�dᣳ[����c��Dq@��2A������P@�O���5fE~t[>�ŽX󇵰;�Ov���q��=�Ħ7_}5�y12��ۜ4ø���tI��"�q��%:��x槟���_ǟ���O�)���;~��A���T�"!&���8���f��{��~����`,׎@íU�v�I�Dkkk��;�CCChnnFCC������������Ѱ�����O����@ �V���TTT ""bR9���	Z��"�Gp�Á��j���L�
�d�`4���e���%�ph�N�NDj\4n���q�ͿحM;�7~z'Rb������A
w����˓�?�ж���'���_>�׬hگ�y����5.~ƀp�W���7S��4��q�?��!3�_N�<&#����7Sb��� p��
g���:#w�袤_��H�S�2!P��@[�e�d"33����-���������b�(((�^�GSS���B��
��v��)+��������ϣ��f�4M����x�O��T*孰�r�8����hhh MӰX,��t���������c�p:q��f�:�!C�w�b����tc�J����q.�Z�
����?��;�g;A7GĲ�H�?�t��p���xs����0+�	ٸ��J� �����I�v��	���鹸Ю��� =U�ь��'
���,�@ ��`��� AP(HJJBAA�긃�gϞŴi����h���cƌ���B}}=���8�3�HMMŽ���i�Z��?>�NgP�:$''��i���J���ꚔY�m�n$��EC�V��uB!���98x��s nmⱙv�̆B̒��\� �{B]��@�� Oc`uX[+�#%�	u �,��A�'�
/��v�8����hA(��Y�\c�1mP*#��1����@ ��|2E�[��V��|cc#�j5���PYY�KKK�L&h��ꐛ��1�����w% "##�|�rDGG���?�0X�l`�ٰg�N��w�D�1��ŝN$��^
+G \�x����vAІ�`����u"p��&�u$65
qW~x-�|�$��~�¦�ڴ�<׆	w!���Ķ��*0��ȁ!���D�J��g�E/'�`VV�V+�v;(�BLL�r9zz���b��b��n��ɞ���`�����l8����*mƌ�R`�X���2?�D"�-�܂�>��d(�����`jQ6,VdR1�N'/C��5�5�		����f��tz��k6�hB!��36'��kD�7s�U �������P��;��B4��S8n���ׅuN0�8Ո��T��
�5��d��$.��f#99���I���ր禥�!>~��aٲKe��!h}Btt4"""<�
�5 @�Pq˜�<y:���z+����X,�Z�FLL���իW#&fr,���Iх�l�f�o�@V�f�'yr v�����O곰 ��	�g"�<���h<�M>:'B���%A�:<,��T'J�h8T��F	���`���p8\8{.� �llݺS�NEbb"d2�'C�f���&8ttt���)�7Q\\<�ބ����z�9sqqq���S��Z��7�a`P�������S�����05�F̸	�a�d܏�P8�'����栁�ڄ��m��I)e ��خ-�! d�ǂ�'N{�����"(��B���'|�GDD��dYZ����hii�m�k􉎎������L���L�2��!b �;�p#A!AJ2��K.Xd�D��v_4	��Y��E����S;��:��Ͱ�]v{xˀ+���=�8���0�GpA,��;�D������A�4�o�ppm޼yB�ݛ������D$%%yҊ�J?233�z�j϶��N���"&&ƣn�W�3���� #-��h�ϯ:?���2�7X4���*�Z >>+W�ĦM�`��!� ��QXX�ӧOs�3�x��٘:u*������~��ף��A�	�O�Frr�ǳ�i���HJJ�08r��F' 8~�8g+2˲!ˍ�R)��Ґ��r]�3�;�0ͽf�$"DDpG��Ek�0L6�PDN>���BTT-Z��۷��>Ú5k&=������r��p��p�n��������|P���f�n����9,n�Q\\�������D�Zy\�יЭ� >F��xn�	 Eg�6��nc�6��mx(g9i�� v�;lE=�v:poZJr9jG/mmm����������;�8t����=K���DO���j��T��h4��8B�7&
�\�������b7�^��;N�a�HX� ��rY;����|=X�ŗi�ى����  ��뚣��T�Tg�B����:P��H4����T*������L c�>>(--���BMMM�csrr<�����P��P�T!�F'��((�Bzz:��󑘘r����p�Ο?��������ǐ	��OXґ�ԁi^�Ȱތ-�i�C�u|]�{4ĈY'��W�PJYD�s�^�q���~�g��#F�^ĩ�f��a�}�CHK�\��p`˖-�?>bcc���ū� ���a��y�F4�x����<���4J,ˢ�����hnn�����l�z���y}�0Å���j )�Aq<���1Z4�c�u�jH�xdB����L'f�����T�e,rUc�KǺ(lo�񕀀uB!�͑+�v����,e���,�~�m�g�ٌ;����B,C$A `���0��A�B}}}��z���7�L&�L&���l6T*�7�K���^J�F��ӻp5:+'Uw�L9�rXymzo<����#׉�X���L�G�(���2��&��N� ����@-e�����-���T�*���␈(�N���v��d#>F��]���� ��� �4>�JP{�;{)�8/���ɡ>�H$X�j `����#�n����P�M�:���A��N��N711����ĸSVV���2�>}mmmX�|9RRRx_kƌ�2eJ��i�2������.��L52;����.�#����R41(n�B�#�wV���,�
����5������F�LK/�8�WC WI��b'���cS&��u"WI��ZQ��:�1����L�_US(�E��i�����^6����_܋{���ǒ�-.��X 0�x���8��=�;Q�ek��ũxv�	���`�A!/�Ei��q �$����o޼A��;��������6(��5OKK��d�*�zfff44M���MMMhoo�.9� ��H�mE��B�����J�Ӄ7�p���uR��57M�Y� 0d�`�:|o�L ����#/o���v�ϗ=6I�U���ā���pq���#����
�4߱q���]����[@��c��]���U���7�ԣ�?��'`#�mS$(��UFG`e�ߙ�����Bt8���Dee����(L&X�M�0�L!�&n����\�Z�
2�4M�_�eq��|��رcZ[[�V��E�i�??�g$d�&��j0+����8C�?>��:����/�L|o�L���8�~���I��    IDAT��WCͳ{1B���i�72����.L�dI�� �C�U=@;�+��f�:<l%9���h%<��h��?ه��D|g�4�2(k��A�~om=�T�� z��
.����hll����bq�b&�7o�k �̅������&Ƚ���� L�>��~;


x�-ߨH��Ix�����{X��g�����($Bb������"�ߧ�H�Ok�=�z�u��d��ɭ�47�����ol i��}��/Dϫ���'������QԞ������ߒ��-���}g/`��Z��CK�Ѿj^�q�Dd<�N�0�r�A`ժU`Y�ׯ:�-Z�V���:O0-77b�uuugԹs�"&&������`ڴi8v��x�0شirss�����]��QWW�)S�p���j̟?�f�Bkk+����6m]k�ر��R��l@\j *k���O���
ߋQ,f���M��s�K�~^Ĩ��z*);�u*#��YS�@�����_7A�"I���"�oI�K��������?����1�\k�r��w����oIx��R �\"BBL$~�r6��h�vU�]SDo�,���j̟?EEE8w.0�J�Bff&����{�n0�F�I͍/r� $$$��;��֭[100 �L���D,Y�}�Q��LOOGZZ���21�B]]���V���������P(��GGG��҂��Fu��ځ|��	�/L.���{߈	���7㙿oE�΀��r  ��]sa�;1�CL%_�@�����Z�ҫ�߾�WzV���|�H����'MTKcc��'��g�#ε~�N�4��B�şΊ�e���6� R�6~��0x�o[  wΞ���� `��q���`���#db��&�nw������Y%	��.�m�@�Y�@D�ځ��4̙3�BWW��Ґ����!
�d�lڴ	]]]hooGzz:"##C����j���a``�glwv����HKKCAA���\.GII	�M��1�[�ZC.�"-%�����S�����w�������]�x�%���U�Q���￼! ��7R��3;�VF�	tΆ?�mP�ꉷce���ۣ�,"/�u?c���r�8�/�"�24�������L���u�`�O��%6k�X8v���N�d.H%"̜Q��>#�29f�E���ư�!�D�@���V+L&
a4QSS���T^)���j���`ٲeزe�G�`�b
Ⴆi������
���-�iu{6			�e������'��H$`��/�#$�1==}(Q(-�D�Nm?|z��{th���ϼ��6T֠��߲N!���ͤ������$�|� (�!��k�7eƥ��?�V��AJ�CH8�+M���Q�.�]�
5D"WH��f�a�֭�����4��{�bժU�5k233�R�8Չƣ��r���ٸ���=�|�X��b� F��N�©S�������ldee]F�F�L]0H�R�X�.�[�n�*�ER�}�F��m5ې�Vf0oJ����N�5��<~?���}���nЯ�|���g�eB�o=`��睋�����:��<5[�R)1<bA(��W.o�0o��@0�Lؽ{7�.]�����w�e̕���F�������A������W�
P��B����ѣHJJBjj*RSS�t(
�RiPc�V�r-o��V�ܹ�78��6���a4YA��=���x�'w@��2���F��89]q�c��k�������z!t��$X��jd��W|� 2N��}.��.ch�ufn�'���}�I����;���`������Ab���͎����S��z�ٳg=.}oo/6l؀��d������\�pV�.��v�BTTh�9�
�/_�[;y�$L&���a�ZQYYT����������G�t@��p8����J���Đ,nP�c�1���3g���\.�{uP��͎X�\��˔�x���;��L3���WoQ@�x�G+��g��M�x+��8�=��By����
�sx�و�(Ǐ�o7�	l!���F�w�D�8��B5���/�8��?f~��/x��/� (r���Vҹ��c"1�#��� �{93�m:��=�
Q2IHc  u �>Ԥ� �^�v�_|�E�cQPP �\�=tww�б���h4
�hoo ��D���C ��$�,�� �˱t�R|��Ǽfڌ�O��� MӨ��ży�Y쒒h�Ztv^Y����ZA�<s�TQP$~�vz��'�7�G���rYHcШ��b�WpT����|�ɷ>~�U�A�����%��ce�_#Nݠ��g���v�����H�H�6t��#.�� $�d�м�����@Gx�7,/�%H%B��xA���47�eY477c�̙���
*�ZRR���rlٲj��f�p�u߾}�繻m6���E||<�V+�9�H��s�eY;v)))HJJ�͎|��H�B�'.P__�L���R�cn��&lذ���.(��X<�)R»����NǺ����q	)���~���ǿ�?JU��eB�(-�63R�dX�`������Z
7��H��w��"Q\ �`�i q���p%���]S�E��ls��, EQՅ���1::
���)e��tP�TA�@܄�|�x��	��*,,���DMM���xӐ]c�����b׮]��SUU�j��³L&�̙3q�С	ݧ0/�k����M�R�Yd��(R���C]�H� ���ƀ��Y�����K���gE���[E�����G_�5�Eq����܅=\��d8r����`�X0w�\TVV�h(p���mmm���G~~>Ο?�۳�X,��ʂ�l�D"�J�˲X�h�G��o6�J���T,^�Ea�ҥؼy3�����,8�իW��\����w��j�u�=��ς���ux�?*��Q
�A��ė��P@?�`'�*�?�	��� �x�Z���D �9ӌ_���3��~Ԋ� ╣V'B�N���-�b�!���?X��bAII	"""<�|kd2����U~��W�r�(..������)�,�af���Y��ƶm�&���m�RRR<�  D"/^��7��p�j���ѣ��[<����R�޽{R��a��-� H��eY�m���H]{�w{���A����";�a�ě�I|P#��XB���I�v\�۲�H��ʬ1,p��¶Q����T�f�	��4$AӨÃ�┾��a���~MKPC���Z�����\.�4�x���bΜ9(++0F<.O��� ���q��c�Ν!g���*��rddd�n����f�����Z�8u�O�; �dZ255�/����
��mnnFQQ���ezz:bbb���Eu� >툃q�ݘ_���~�M�u�0��ױ9]��nB� �WOHpW�y��s���W��'Nn�U~� ��v%	�T4T2Bf'�a+�F�j-	���q���j�=3��n��~�F���LO���g-��cPA�5_t�,�V[[�Ʉ��X�V�;wÄ���ގcǎaɒ%��s�Π<�4McϞ=�(��;w��u���#G� 22�'. ��Y=�S��|�r�~� �����G�N��C#�Xמ'16<��m:����H�$Tc���aK�����	�}F��(��i�((�,�F;�3�:��Z
�ɠ=sCg%���Ğ��C����qt
��LJ��?�����>$O�w �Jq����_SS�cǎ�o�٠����,d2,K�YNN���:�ܽ���HLL�ʕ+��'�����X�V?~ܧ�g�̙��d8y��U�S���Rttt`hh,�b���X�z��"A�1c�o� ���^��	���������I9�c���]x���2��4[{��br<��A��D���'����"H��c���ܳ��2�H�`Yv��ӧOǝwމ��rTTT���Fvvv��4�g����$&&�$橐$���4�u�]>}J�yyy!��W
���1c/^�)Y��l�3|JJ���w�P�!�Hx�1�$ s�x�1��>7U: ̐uB,��C�)�@]#;�y��bB���j�N���`��S���h�p�BlݺCCCA��)S���i���C("55���hii	zϚ�ছnBcc�_-� �H$�ҥK�q�F�L&���Z�FTT�"��p�j4�L&���]�x+D)
TTT��� ��҂��"O����������S��Frr2z{{'�7e����c��dp$��,۷o&39�̓�f���	�bH���X4ݿC0+U�����C3-Dn�˦Oޏ�F�^� @�4�@bbbȗ�l6����S\t�=��R4����N���j��n�j�d2!22ғ�;y�$X�Eii)d2ل��R���ŋ}*�1������~_NN��������������3���c`2�022�^5��p 	�r���D�#���=�;�$I<:[�mg��hQB��կnc�p	�X7% �g�"?�����~�pxT�~�sWW�M��e!����Q̟?���8s�L�s���QQQ�F�$1::�s��%S����1�|(�J,[�UUU�hƾÉp9*�J�~�������!�˱y�f�u�����y�9�X\���{���3g���B���m�1�[&����n*���d21Vύ�Xt��6a/z�")
�*)
& ۿl6����Ijkky#++E!77��u�������g.(
�\�III�<�\.��ٳ��t��p`�޽�i			X�b4h��PZ��o���V�1m�4�m�����~ESiii>�\)Wo	����Z�N���H���r&���g �X�N�QO#I�˄Ĳ@��@U� G{(8�/�r�s:��i�\�AM.��!�J�s�N�L��f�.T
����χP(��� ����t:��S������ռ"�ؽ{7.\�H��Q7 �������*�������O@S  ..�#���|� ���AGG �I�Lƛ�d�lC��.^�r�w��(B�E,nN�1-��8�S�.�)�pv�
�`���)t : cA �
�
'nJw�:���n���O�\S���T����eY���A�բ���S:��x��o߾ݳomm�X,F^^�ry@��'N@$y<���N|��GP�T0�L*$�k��Tl\\����V��c��f��Zvy��\$2�����яW���4�8'|�D0/Ņ�r�(���1��\%�F���
j*�\�v�3h�7b�,~8ݎ�E8�ͿI)#A���oH��߶�SV��R�"!F�%�Ů]� �R�F������@ ���6�_�f�_�͍��Alܸ�sA`Y.�w�y'�v;v���Y2+���AHJJB||<�b1�V+�F�k�Õd�r�f7�fxov�ߘ/O_�(�6�6����db!�߃K������=�~`U�s��{#)
OT���Y1ZG�ߏ�� OE�e� 	�[�b����g%�iYh���Ϭ[af<�24H����d@Q,��h�b���J>��@zzz��� �e�P( ��������(++CDD�Arr2rrr��䃔$K$,_��s6��lصkWX\�@hj7�������͸t(��\MS�)�JQ$fW��d!R���G{Gh�8Eb�l/�.h�
|{�Tt��h��}h��Qy����,���!ߛf�k'$�Yxv-J��S�7n �3Ŏ?���3�����ʏV�ݧW��ol�W����\ I��qhj㖋S+���F���Baɒ%�(
'N�����=hh[�l��hI	n2�P]]���|H�R�9s���A�iii�ԩS=�8�������A��3g��3À$IH$,\��֭�x��Ϸ�l��@.����q�V���d�&�1=5z�C�c˨�::Bz�E�	����������/=��Ƭ'���)�F1X�1q#'ߙ��'��/Ω{A���_�� g���=�kvw!�����l?y��nQ&f��cXN<���l��[�ݍ�%���ƃ |�#���U�\��j���ctt�f�����J��I3��nGCCFGG=MO�:Q]]������`pp###8t萧X'���a4��'���>�P��]�.\�\.�������0�۳g�� ��7�sKr�
������=�`[�]�̲��~�/����e���y|��> <�ʧ(��+�|��e;9�L�9�-�bW�䖽-Dve���M�T��J�f8���<� f&�蠁��l|�՗�6����3�?0+������~fjhlk�E�bs���+���V����C�i��!����pҐJ)44LL�8�/ߙ3g�p�Btvvbǎ��dA{��r�������C*�bɒ%P��A+� pr���ׇ��H$BOO�'���ߏ3f�������CVVքRr������ӵZ-jkk��Ϙ1��<�V�YN�$驁��w
t<��n������./�X,�D,@O� onͷ�Ǩ͎�?���j-vf�l�#a����y����S7o�Uo� ���/�zg����xR�D�v��;�3I�'�IU�g�!��×^�P���MO`���)f�ń�D�6�>�����x��J���q~�M]P(� 	14l�"�oぁ�BQLL�v�'�###P�T�?�e4����`��M��~�i����Krɒ%p�\��� ˲���nA�|�Ɩ-[�d�N����_}��_�5--���~�{�$&&�)�v����^��ma�Ӆ���RF�jux����}��:��!����c6��=�緿��a�}��+?P���-Y1L���\!�����XAF�z�EO{�Q��	���;>�+c���U;bB�~v/m�Å￼�<�m��;��b��f�x�C�K^.t:\.�Ν�ٶt�R��SRRB��UUU���Gdd$���QUU�3f�f�M;J�Ҁ�-�PSS���5566z<����	`��X�~=rrr����H�^���O��xtuu����m���>��EEE��yݎ_��]���f008�� �|��/��6��O����'�����+vް�z)̛�ۄ$%b��1�^��I����g���������S.d}��T(��@��o�m�9\��օ<��GC��.���~�����l6�ݻӧO�L��!�4X�n(����_}�U���ԓ����Dh4���{R��<���8��偢(tww����`Ϟ=hk������h0��0ػw/n��f����1G����q ����=������&�˔�����{k���Ä/ydf��i����6�{Dp�ތvҀt�
���:/���\��	��%��eT��
h_xa�@L�~׳s\�b� ����HT��x��ڱv_�:}�BvY���������� �j5�Zm�R_K�,�|����?p�׽!�c��@c�����ѐH$�����d
K�y2�0����Á��.OAI�>��:��'�8����p�����x��"RgE⩻�##�?0[�܍\�iαI�!gA�U����6n����0BȖ�]�2�;�%�'��?��	W$��ݍ�E81�$4B"����21��|�\�B���z$����<U����111~EGWC�h���(..�IǱ,���6:t�W��d�eY>�쭨��Z��;�;x�V����mmmWTl7P$�W|n���c��>	�P���o��2��遐��R;�ș�E?yz֞�}9��	���ocY���g��$�����j��~��[���������eE�~?~��&Ц=�.)�ŭ%����c���~������p��Sh��rL����H���ԱZ-�k�`f��bUi$"��U���`��M� �F���",\�&�	;	�9⩢��d����e ��;��� �T�7g�TTT  >���Ģ�"̜9�o;A��̄H$¶m�B��^p7�5��I�Faa�_k30VG��j���X�\#    IDAT����X��J���v ;�?�98<��k�hwh8s��ұ�� �xg+'�s���w��'k���y�Ĳqqc	��M#�>�R���~���}va�ʶ���3��:C4�(���q2Vx��ޠz���l|������{��o�*�����!�K����!���C�� ��2C��t�Ot��7��`g����Rp�ƞ
�q-[(���N.�˓��*ccc9�a��,Q$	h�FNNNHw]$�E�������r�p��i��vL�>:����(**Brr2
E�b)`� ��(��O}�8���QRR�R	�˅��N�8q�׵].X����g>JHH������l�t�Ŏ��Eb�b�{7�w��xZ>�8������ۧEfc�/VN�m����?[9"��zz��'����)Jڕ��'���櫞/�����b��?D���U�ߏ�qW� E��l�9+�ȝ������2;a�A���8�v��W�.�ޙ�U���#�����;� ^=�8��w�u���3g�����b�
�e�z���֠�#�fለ��������g1s�L�ٳ��-
�����t���hrrr|h�233�����?�<�r���	v��-EQ`Y����=p�d�QUU�C��}�����g��X�e.t�1̦\������U�5�����:>+G���c'KXc�L�B��|�Lv��x�>��N�q��j+RA�#*;�/0��,�SK�$+��hn�����a�֔n�����0A	M�
�
����������H���vOM����EQP*��e�L�H$�	~zG��̙�y�D"AEE���$:::�}�v,]�'N�@Wץx��ٳ}�L��X�D�μ�N�f�ǿ�naIF8jr��c�:�K�LC";���%	 1��l���6�rz����B�E�(��΅�-T[��Gy釁2l�����,���h���h���!tH��V�͆�[�[w'''#++�Wd~�������b�{�P�TA������|���b۶m���BQQ�����lkkôi�|fm�N�A3��
v�����) ���	j333q��^�½�����|<���lL�2��8�˅�Ǐ���FA�k��k�+`iLK�]�e%E#��(�,̣3���,~�p`�Y���)8��>8+���v�9j�Baw�g���πƀa���E�+߉�atH�`SSp���8Xۆ�G_
�:cs8awr&K#Wԇ{f�S��&�hmŁal#CЏ5%�I�cY�'p��������d��Şw.33�w L�VcŊ~� �PUU�X���\���>8p v�---�����5y�(�wI���ƹs�p��73����Ec�ARR��:�8z�(��("��~��5K1����2C��x_^E�X��O5`C�=�G��tK
}	BA���������^;!�C�ds�'s�f�MMB�
�t��gX��!j�n�q"�C�Ս���B\�+
�	���ӥC�W^�,*�` ���`ry�R)��^��|z~1�/��`@?rss�R�x�8�\.TVV�СCW7�<���l��(�J�t M�ؽ{7
=݉��$�g�������MX�*�RUx.p�F!� p�&%D���TC'>�N�<�bw��ˁ�I�*1�44�d��
 �Ȱ��
�Z��m����k!��	1�R��B���Vl"1tՔ��Z�X���0��t~\�\O{f4y��n��˅���v.7f���K$H�RX�V�T_ss�'ة�j=� �[0�,�m۶aŊ�x������(��3�5x�Y ��(Ti)$E��Q҈3	����@� ?5% Lv�a+���������:��Äd�X���oO�܉Ҟ�\.�'p��!�4}�l���`0��px<��B��z�]�����B&�5`�X�y�f�v�m��ؾ}{ؕ�\�i��!�c�<��������16Y�ƠJ��ۮ)��Ƒ#G|>_���D��,���=�?))�O����߇��{ip9�n�c۶m�D�֦\�O>��	�?Ɓ����,C�X�jސGH�RF��(]�7����^�w2 �X�D;#ݰ��}�pA��*""&�z�z���G^N2Ԫ�4
%��M_��7t:N�8�O�FGG�O�J���&*�v� P�UQ���X �V�m�S�_7�pƀ�H$ī�ta��=�"bG�����13�Պ�3gB �eY477�11�F�[w��j�ꗋ��x�X1<2�F�ˉGk���2o_m�eT�K�� ��.ftdP>�k
����.MMM!ۧ�N��^\�KN�c(�Q2�l��N�et$F��M�Q2�-ۉ� u��Z�h��F����"3]���HD��
p ~�/�w�c��ȤB��tv^{��$�2��YN�9bX�np��`�|u	ܕǏ�=5�����8�Ma�y&�D	(H�B�Z��D�D��Vx�^�j�!	�כ�:�|.�\4��Ct�6���Ӑ��!���9��ѣ�� ���(T���0hi@�=$|�؎���F��dJ��T��*I.JO����1r)Z��x��-x�G+����>��⺰�d�f�h�|�o6���ȵ�u�E,+w@��	�*p"R�b���`e�3lC�F����'�h�׬�������Eϐ/�k7~s�Bl���7l���m��kn�����]�� .���;f"R:����}���W����ɱX��l�総 G���*I �g��(Å~3�3Z�-̉����-���ĨL����3�:?ͅS}zL�cӳ-�b�o�E�#�V|��<��/q����~x;Ԋh9,�����@���JX�1�wF�B��	��xp~ G��`�f&��`i��@��4;h�-AT�؟�� �;��`Ł �3\�q�a;;@=���W?to���g�ʉq|��d}�8	 K�\x��� ��6���3Yݟ���� gqOҍ:R�8Lܵ���<}�=��o����)b}܀H���N|����M�"
(Ps�	��oC  �z�M�#��A3�ל��d�E{�q�5y^a: `��1��yS�>�)L˲p���ߟ��8T�P��w���wށQ����Ζlz)$!$�л�"�Q���Y�<O��]�N������SPQ�r��5��FBz�dwgg��ǆ%��$����;m���|�}��y���)�Ue��=��1��8����݆��{U9�P�H����-���۸�A�N�lx�!n������9�Y�>}��O�c�KS���8or�B��R�u')�&��9o��gF�x���9��/��^���P�������3V��J��F�{���ce��n7�*�a�/��q�!�����q<^�-�O���9�<{�H��^�f��_����#��),��i���Wƻ�:�Ӗ�GKJR��N�j�h�C��_e�Vw�#��5���d��`!����g]�+O��}�XLh _=?�CfݞLb����Y�_?�����>3	?C��޼
�-���`�3W.W4��bnPO�C�-���8���rS�~H�@a>��2�ZȜ��QTa�__��?�߬!����?Y�M���$�&��8�U���ӖԨ�kh�=^BA���
6,uۖy���rL���GLh ��[���_v1�m<��2zv��sT�>���W�,+�ͳ�f=l�݆���^��#?���d�Msg5�q�m�oLsD��J&/���`��?��������Y�a��ZOe-���*���&�gf��U>�>����QՠnAe��˖+-uq��6	�n���v_�~oz�dv�z�Cx1h����pͽ��Y9��F}����1�z�;��Tȴ�H>{�b�=g6�����1MM���d�hK�`���j|��d2q�u��i����I�D,P<z�=:��.]�1dKHj�S�v�S0��Ld��=,�|�u{3���VC{8ݕ�����%�lTCq�}���湻��y�AQ��T�N��(��i�Mu��K��H����|~2�Z��d��>��'o��'nc�+�\_bC
&���:W��ĺ2��/=�&w+G���I������k�Մ�"��#@Ld7�d��dg$�P�I�d��M��f&%�1?�V��"���dٖ��q���z�{Q�^dh��|�l3��P�S�f�z&���G�xf��o���y����B��m��������	�A��Qe�<���wfzT|���ǧ�GI�6�^i������t�Ld�?7�}م�&%յ6^�:���y�$g�+%Q�اE�2���"�,v�c�1�{V�^�����VX��a�>��#��.�K��N�T�OP`�����E�#��/��(M��/9d�����n���H���+�W��b���-��J�����a����%��Z���?���a��,��h�\�U�-y"�tq�D�k����tRQ���jrl�S��~�'zD8.kX�`s�ާ��>�7_y��fҐc�͈M8+D���!X,�͛�*O��q�$�����I�%��H��b�1D
P�}��y�K��f��V�p��n�wq��*�J�~�y��%յ�-��Y��8�S��TZ�ë����B^�3Ve�4A&��ԃAT�#$�/�[Tv[Na�Vg�^;�|����9s�w344��䈁��GR`��x�&���H�4��E��(VI��#�`��y�>*0o����j��-�(k}�K�x�ß쭯^\mi���F�������O[}��Ҽ[��%��:V50�k+e%��������z��[��-E�o��_仯���y��u��B%�5,ڰ��*��5(5mS@C���nwPT��ߐ�,yV>K�<�'Ȥ���8���FJ���d�Ӧ<�R����턙���Y��kl�����������q���7:Y%pS������
s�4.�����R����%	2�:9���E3Ur�tl�ِ���PvR�;�-���;3�s������������?�ᣍ�3yEo��WT\ɶ�G�<��}1}sų�$V�m�����DF�^E��5����uO��Kr���ٺ��g��?�5WϮ�+�d��8<j/:T8V�cC���"�ѵ;����P`]�Ⱥl� �J��*5�[��.TztK`��||Qqe�b�)&��c�W)����6-~�]/cof�bp��C
���Qy��Y1���t�{$������7)�z&1�����oHΉ�'��/=�g�=�~*�~*F�J�$PZ��X��-vG�H	�Ws�s���T[l��H���J`��͊�Z,6���N����.�dj�Y"�,c�9�o��oEQ�Դ���B��*Pnm�oGa���p@��{N�C~,V�U��5���)Q��ޡ��
��0L��1�'����$_((��]�JzU�Ҡ,�_ҩ�"SSc�����!�n�厡��ͭ��(���M�l�Nā�D]w���2��X��$�N�c�	��;�U����� �0K���d�(��d�u��r!�O�vj�*�*��9��(�9���&�+L�HVI����*sv��U���D�V��f���n_�z[%��xTA@A`��3��>1k��~�N�Q�h6[����3K���v�)Ne�2�`�,��ѫ��U^m����yU��F��]�ΝW��_J럒mMF���֎��9��έ��kWU؝�:w�j
Ϭ���4��*�l�<�כֿn6 �{�={ yj%e���ȓ=�R+�s8W�$m	�#�?��'��l�A/�)���}�X��:��e��$�!���~�U;����;��8{O��?���7l�5ȫ�E�x�h�3m�����O
	4���9��&�9<�.�R����Sl%����g����\�Y��S�(�>���ts ���s���MƠ ��5�(bD:�;M��ʖ�M�a���8CT{kc�����>�l��t���UHM��'E�������H��5O�49Eu_��2��s,��#Fx~�
fY�]"�Ut��!nV	0�X$��Z�%";D�|X�荛����O����Y�q>z�z$�лY��o��F�]�Πi�4�v��q����7Z&5\!Ĥ�W��	���W�cg��쌟Y���M�7�ܔ�`H��#1ĤbRIU�.EbK��%��X�������<\�qU56V�8�x�n9��-i/b���54:1
�K� ��*af��{L�ĪL?g�,nԤ��L`'��v� ����+|��H~u�{	B]Wt�փT֜^��F3m�?��q���o0�+�*?n?��J��H�R�m�O��&Fw�H����HM#�F� Ĥ�� �Wߵ��0+<8��ۛ���X�5��YQx������[\��5���OGP\i�\[P�q���ſ���! ���]�I^��R���gC�dj��m������ݫ�����)*w�����䓟���'x꣥�~�~�u�E���=s�H"�����/�6����q>�q<��S^�؞ɧO�΢��׿�@N�O�4�Li��"!Xelw�o�{&���z�S2��qP��坽�x��p��KV��sQ�P��� ��	\��Jq�@~�o���م,�z�m�sqԳ6�u,�y�w�d��q�PZU�򭇸��^Lٟ/مMj�awS���b��b��2ݏ9��ueV��o �$z�$)�.�b{U��3��}Zls�~����#�f��FN��O�.[�?F����#�d��7���g�3vX:��Ai��v�����5B�иI�#*$�GO��7�q��H��/���Ϝ�p�퓞x"2)ر=%Tv���	pE�����g�zܩaf��@����B��G�μ�Ί��Ow�����#��E(=��R7���6ݧ������.{��A���|J�2��8߉	��`h��(���v�cʌH��W����{�ho��/�?�n����w��d���jat��u�+J���7��$)^���Jx��옫�)D������
��M�<ݗE����07��9�����-�}����f@�8�{���6���7�S�c�7!�sxP-��sLn��>{���s�����o6A��궰�C����{�$�C���M5���6�~c��ohP��Ǖ56	|)d�~����7���O��Mj��L�vf��L}�kL��CV�%�X����^��j���G&�/�]��kF���޽>�/�uZ��^G�� ����r(�#:�htht:����;� �7��O
zQǨ��>Q̡���T��K��Du`Ёg:{��bPᵢ��x�b���N}����c<P��z�4��8NK�i�r(��3��ve��F;qy�df?qC�E�M⳧ng`�� ����X�/��kUZ=������N}<|��jĨ���^����!9�:T�3�[��M�O����^ϑ~�'��*�7?�xy�d�>3��u{3�:cV�]44�7N���u:^�z�������*��y��	���[����(����T��*/j�*�W�oh��ل�M
q��p{�U��ތT�r*u$����="�O���>m��M�N�QF�;ݯO\��]�e�b'��|�l9��f}���Ɋ��]G5!��ą�r�a~ݗ����w����I�����"���GIz���f̼�z��}&�s�uK���a��ǋ'�ט��,=w��\O?���;ɪ+��#�m�p��@RBP��0������"*6Ifٖ���G\x��P\Y�%=5 ��̓^ˮih\Hd�1�W2f������e�5GϕI�G� W$9&��c�ͅq��Rl6�#9����A���
�����B�ce:R�d:��)�p?�C�j��r�����2����|�hA ����[��oQa�2��/�8����44�'��M|��V�]��7c�w��3�yhܥX%eվ�Ѭ<�g`�L��Y�� �?>�qus�X����˺!�zU�Ow}��{����6��3�{g^�w4�f0��و����0���l�g?$���Ϟ��62���8W���  �IDATJ������~���:SG�OG0(-��3P�OG�$��Nc�K/Yz������m51���� ߣ��4z��h���A��_�����'+���#��W� xg�z>xd"��~Zj��ź=�y��𫗁�ST��+�����)�"�B�G;���׎����E>�c�����d�AI��ۛ��U���T�S8gQ��G��0�w ���{3��"�v�̷��xݗ[\���.����M�􉒛���H?ӳ>G��R�.�M:�9`�A�d��#�3B&�O%��vgI���"b����N#�G�_�?���5�Y�qp&iL�~56�jk�LB54:"%�:��2��'F!5�yo�Ξ}�E`_�HF���c>Q)�
��ҳ&��uW�e��L^���go���Gr]vg /LE��NL����Z��ZC�!y�:�u�hyM$7���n%�-�Ȟ�22���g����?og_va;�LC��@��lE�[M����=�=���-o[CC��Е)~hY8SCC�Ca��w��=/�RTuFz�M�kh\d���^&'h��(�Tt<���?5�444�:��n�f
�nW^ ��9n���F;�����麠��7"/�2��ICC��9K(h�3��*� 7��<������SxA�U6jhtZ������X����*���Җ����8��qw?��i��o�
Oqm�&�v����#��X~�
��h����q������O�#�Lk��jhh�]|�����m}M��O����7�и 9o�0_���R	6)��A��۪����>�S�+��J|�B�Q Tt:�,Pmȫ�5j��q~���y��ק:0x����Գ萁�v��4�pS�İxQ�z8�:���Ve�ϰ��ƹF�vfBw�+�6���`p����Y[��E�ʃ���ub�ÍiqA
s�}v��h�>f��3�#d!����8���YU��P߭}�ק8<������۲ض+K��?�N2;i��.$��A;2����b��|�$��j+ ��}uO�C]����C�sCupI�{�ς�*~X���.����f\?�ͧ�k�,�-_��](h=�v$!ؽ},��%�,f�{_��1�b�m�;¬bn��s�K �6��f%)ڊ�M��A�M�bj�m���a��N���V�Mڑ�j�Z�]:�c�s_��-�����s��V�����#-ƭp�A/���vL����i��h�vd�	�����f�����a��<�6�]"IJs;gO�H��܊�$l��p:Ƒפs�h!�H�W��t�}^�����������#'|���d �S8{�
ڢynt��$�����3��+�G��[��Ġ�(ٞ/20�� �>����˭�h�e����D׫�B|�����E6����?�gxzr��|�t/�s��
��c�3w�'�W<�>9E�m�Jg��/��w���K��Z�ѡ,���|�t��V��hbЎ�*��k��VbT��^l�S}�Xd�~C�
ڶ%�xw��[zJ�:T�5[ϒ#�&�����&U�%���3�;�q��5%��~|�������7c���z� �/�2���V\K�vFQ�ǣ~�4�&i�AEP��*�]!PR����$��n#�~*��
��*:*�(�ёY�k�,ɆȲ�+�?!���W�M�1è�ٙ�p��1���_J,6Ɂ������!��{&�$��@r�<�C����,�}!Pn(�^mm���*n��\V�� /��!��������K�>�_�������f,�Љ3�v$��g}��þ�BN����v$��
�͎Р�y���M{�rө�g��vi�8��-]��[B��t�>���h���u���O�j��@3�M��@?#�
�-X��}Y<��G���Rk;=�z��q�t
`���,X�۵/!2���I��ۓU�_>��nhaЋ�?�fbBx{�z~�~�E����A�(�+�$�(��
l���K��$kyj�+�"���߮�Y ��#��g6IF/
�7�fV�>ƸK��
	`ʌ.AH�#9&� �Hu��]:18-���Vo�Ш��%��@3��"$��Np^+.<�@���}��51�W�r��w0��^�il7��I��h�R%��8�`���x������uu�v�
�-��_���Oড==��x ��_������Wa�S�m�O0e�|*,V�]��[�E/���jl�=��q|��-(���`�������vT�o=��[}�쟶r4����øK�9�WLnQW��ʬ�s�̯��9D���Ɲ��z�YvzF��d�ӧ�`���t�u<��2l�̵�}H����t_���+}9P:�a}}1�Iv	��:���:Ec4�$�����';=�k�c��z8��;�
�ƴqÑe���%9&����Y���ys����W��ɣ�a�~�e�׉<0f�?u����$F�"+
o|���56���*jm�.X�^�1������j6I&���ǯN�b�5��xyo.�Ȕ7PPVůo=Ā�33��I���������5��Z{�	צ8��
�W ;�y�{]/B���%���%�v��|�[���:����K�yk�Z ������K��x �G��ޕK�K�1���*�&g��=����6�'9��`�F���������W�X�;djm�~g�8Vc��|-�Y�M2���e�e攺� �Rcg����0��X�+|��Z�:G���* ���3�/(����:g�g`�w�j�g�uU�mf[����i,�۽���W�q<ߵo��?���Y��}�T �?��f/w%x�M��^ ^]�k���!��*6p(��9��Ap[�Zߴ�����BߔX����QaΠ_���b%#� ��PRaq;���Rn{y.�]?�N�^�q�e�4�Y� +*�(�JA����F�Ǡ1�"�>i�W�Oe`]!%6�����t�~�K[�[�ihOws�z'�0�^,ڰ��rso�U1�d��E"�bd�C��fD[w�`�d�&GЯ��K�9�@#�w�����z����n�b[���'˼�B���_�pm�v8�W��!-ι��.9=_�ccЋ�zp<!~l<��&׬��2<5uXcs��W�p�Mr-��?4���U��H�z�(�C��W����:ǎ7,6;�u1� ?#���������v�ql;|��d��@\zXO��R�"HI��8f����R�b�����z2ぱ�N���қ�/w�b`j<��<��'K�	��PTK#_�F�B��-0j�C7]�C���p.���۾@��.u�@�� 5.Q<���/�����+ݓy�;_�����t�~����lp-'�ìo��iTU�7������=dUUY�7�5ǘ��<�����;_��,V;�����A��eյ-�j<�bP\���m&��g'�Ͻ�"�K���5��f�����i?�+�y�f�q<S��T�pi/F��vζùL����}�_>7������@�	�y~�r��Q� ?#��{�����ė>%���t;P}�ni�(*�E�+&䍭�s�����X��MÍC{x=g�ǻ�>�S��/|�z�~_���E��_��,u;wO�I�d�l��*��fz�x乴ě�����>M������G�3��v��D�$�(E���
Dʭ�7�ځid��-��܉NaA��q���ueX�D���f��M��	d��0Ꝃ���	~�~p�{�1�z���b���MX��ݕ�]�0����7��J��^޽!�9�����B 0�G"W����,Ov�c�$(�/�31���8��V-jhh �hhhԡ���������#��ų�\s�!s�����8G-�hb�qA�����%&ܧZ��<2~�[FӜS1�	����[�X�
P�R�o��s��A%.H!&@9�JPS��� ������{���s�,G ^�z���B�i��-�`T#�����(�ᐡ�\��� �e	Fuqbr~~E�C%:�?d����:ha~*c�I�9�SmX����L}�l�D��;F���be��>��a���������>|�ʷ�.f���P'�}���*�� �D���<6�FT@���-]bb�%��^zD*<:��Q��B':@�a6�Ŝ�@�����~�����Ldp +��)�3�]��!�Ǜ.�p�j���0�r�(�ݶ���w���u.4κ\��g�s����s�$;2NPV^8=&���LL�eP��и�=�M"��׎��t`r����W������_�?��Ѫ9�J+�v�:G�2�o����4�����g&����y�cy���ZԆ���\t�!���o>���|�$��g��`���t<ň���a~*��μ���@�0����{z#:�.}S�PT��s�?�_��z��lQ�-�����$&���S� B�32g5fjT]]�c�%�W�v�e��{N@b�����x�C'@|�i�����=��;I	a�w�q����+�,��]I��~�X�2K0E�',���5��T�|(�=!���r�k�c��WZ����5
����.s-c��O~����Љb��y끱�$��k����A��G�Xo�������"O�z%	��5)˫�Ǽ�����7_����tӁl��@\D0OL��;�����]����!gUt��O�����o;���:յ�C�d�_����:�D96���}�S_�:Hܤ���w�����^g�(�q��Uh�A�A �l�H^I�ڣ�*{3��o
���>xd�GA��u㙏��p�׶���ځi�2������&\�Zn��G����TwC�у����?���}�E�~x�tw��ط���b��׿k�}�V"�z�S ��Flx_=7�M�N���A�U���?����H���p��Q����b�z����?Ӊ�.!8���E.1��:��u���Q�%�6��̜2һ��~=Q� ��L?D�SRY�u_^i���ғ��̚���ُ8�^�1���X^��71P��?Zʋ��D�M�	���~{�@�Ƴ|�A���*U�K�p���-�u�5|�q�S�n`7jl�6�eDP\ai4��W�?����m�{���*%�w��C��-��i��1���gY*l=�gx�� #F�fǞ��R�D�-�)�V��ek� �U��f 0ԋv)��a^������|f�!S\i!��i�7^�:�����K���ԅ��MC�%�݋�����p@��������m'����7�����J�� l;r��q��n,��ݮ!���{�>���F����n�b�{�E��]�6e�|;�Зu��5�k	��#�G(D����uE���
��:dU%���>>6��� 
���v� п��.���Es�Kl���{ǓWP��1�%�{��Ӌr���DBd���S�"�f@��'y5����d�s�)��Paqw�ޟӶEqTU���g�ƹ�,&,�{��^/����"w^5?��ެ�d��!��bPL��@��㦀:�u���b�t;�#�#�eV��{*��g�p��ꌇ����zq�h!5�v�È�<m�~��c�NT��,(O|lo�Kfv)~~z�u�B_��P+��˷��^��s� �9�g���f
n��C�C�O����$�k�b6���7c�ˎ���
f�w�6����O\D0����jl�����{%3��I�yUf|��A�	L��5��NǠ�ߡ��,���5�;��{�񗤳�X��cZ�9�@���v�	PIQ0�U
�u+�q۶;*p�L�[���E���rGģ���OD���qyU:�%���`�n{S���=�ݞ����y�  n҃A+������Q�kSǠ׸z���\3 ����r� �l´�[Ē��<�S#���1���Ⱦ)���Ꮯvm���|�#��,�����)TUe��?QRY��C\3��G�z~2/L��&]�v�/��q�_���-�����C�:z��1?n?��f~CKi�_�����xo�,���*�:Jk.K�2���8�IK��rˏv��
Uv��`��ffG�9`���4l���/��	�����z�N��g"o�#�!,�z���&�CtX ���y����܉��<«�%�dEe��CD���΀\Nq%K7�d�U��� :4��?ow���=Y��=�q�
K� ."�,SX^M^i�,Z��� ��w���RKay�똙�1�gg��b���CYU-K�`��Lʪk���#��GPQ}�܂�j6�f��l�vk2��->���ǔW�a6�Z�����������m}�����C��e�|��ԡ�g����V��cz~l��]��Čߏus VT��l��5 �M���甜䐙��^�j�˪\�q418G$�(��� 5L� Bi����zVg�u�ߩA�':'��P�x���L�DF��Ⱦ]I����jgծ�n�t�^�J,�ȁ�"J��O7jx��������hhhԡ���������F�hhh �hhh�qڒ�)6UP_de�N0z$��2�i�A��%I���R떒uPl�cٕO�����%��Oo0P�E`��S5���	���7���ӧT�� H��d��L�i�?&��%�4V�3���/P4oP��f]�hÄ3������8��{+X6�&����͸��zg@�]*��SbPXX�$����ш���`�=YP�S;N��y�&�SbP\\Lmmm3Gw\���Z$�M�"�%>44�%������vn�����Y�t�i̘1��n���6UUj�l'�+�/��;  `��(ہ������,7��Ձ1�[�*���2Y�_�o�Vi����@�+��r�0�h-�V��WWW,IҖ����ڻ=�#�6m� �⿿�����ƍ�����@m�ل�E3r��m}�	����l6����揾8E����LA�Z�ʯ��sѣ��L-���#���ŋ��			�<�j4�4h��h�����j�X�����Q�8+bP����*¬�q��UU��L��H�����g�w{�WAP���d������.]���m��YX����gm6��|�OA�Ia �u�ޣ]����(�8v��?�Gs.TF���}��+P����y.��߮�Ug?�#p���w �l�׹D@��r�k�ڻ�������>P�u�����ů}Aݐ�����qs�U�NPtCT���	�9�p�J�}�e��9�s@��'�"w��I{�C����5+fz[�8JY�����    IEND�B`�PK
     T\��  �  /   images/858a2a89-b1fb-4d30-9067-568b89f7eae7.png�PNG

   IHDR    Z   P8�   	pHYs  	�  	�Ǡ��   �eXIfII*            (           V       ^   1    f   i�    {       �	     �	     Pixelmator Pro 3.2.3  �      �    Z      ���  niTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/"
            xmlns:xmp="http://ns.adobe.com/xap/1.0/"
            xmlns:tiff="http://ns.adobe.com/tiff/1.0/">
         <exif:PixelYDimension>346</exif:PixelYDimension>
         <exif:PixelXDimension>259</exif:PixelXDimension>
         <xmp:CreatorTool>Pixelmator Pro 3.2.3</xmp:CreatorTool>
         <xmp:MetadataDate>2022-12-26T23:32:11-06:00</xmp:MetadataDate>
         <tiff:XResolution>640000/10000</tiff:XResolution>
         <tiff:ResolutionUnit>2</tiff:ResolutionUnit>
         <tiff:YResolution>640000/10000</tiff:YResolution>
         <tiff:Orientation>1</tiff:Orientation>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�Z��  �IDATx��]x��>[�齑@	�ATDD@�+^��{U��-���**�ް��� (�{%@z�mS����_ذevwv���}�y��ݝ����~�5u?(�g<�WP[2��e��2��D��P�(�=��A���di�#2�4II7r��.�ɭ�ݯu��-�l#��I�]�Ó9�y��	��_�p_Aa�$(�\vifZ��IP�?ɮ .����
�!��#��g�_�m<�]��$�ت6�J��6�d^S��S����#���K���I�P̵��?��m8R��.A,�f�B�ea��!G!��l�{���'�u��t-��K�q��[��Pȋ�6`2����#�-lu|��ܶ�~x��+>�k�`���0�n�@�_�L'2dx�fOU������˪V�3�k�W:?�������=L��m�/C�׈c���M:��K\���\j8t�� t�C�Hп�H`ɐ!���a���-Mw(f>0���'����Bg/�a�2,���MLÇ�QO�G��F�5�~;�R����I]�_�溺#~=��Ӱ!]����v7;QBg�tAI?�]��&�aa�O�K�ud��Aج�	�F��M��E��RO��o���xJ��K�����~?fR��.��weSw���Si4��|`�����"l���|�=֐2��LK�>dփ�7��-�]�;s�N�A�e��	§�@��<2�L��M�����{���u�B�|$��h��=<��2����k��qd$SXhGf4UV7Pn^Y��@C�PW�_�32��%�M�V:�'�ĸ�ta���/�z�WO�r �� ⊇S�F�O��YuŬX������{��#��cE��G�t�������m��w�/�6$�tZ�J�W��+V��Xg�]?HmVm���K�~⨷o���.{8�l��'I��	)d6�\�xr�WO��^�AȕK���{�P&2�'bf�ꈙ�ϭ���|�o�"�>n4
?2��?ɐ!�;#ɬT���IM��UHy�t2}��(|���$C����FZE3�O�R�$�B��G�p>ɐ!�,�bb�J��&���^)�Bg?0���!CF�����YK~k�v�*w��H���ߛ���\r(C�Y
&����g/�[��2��tOd�P�Uﰿ�$C���A��{���%��K�����ɐ!�'`JȥK�o�n��bO�$���Ì
��H�=
��ȩ� �5�%�T��؟^$C����S�������O��A����˝$C���%��d|y�7����%�`y����
2dt��"�h��n'2�da�@tɐ!��B�
�r�mS���@��<���H�=O�0(�c�b�gO���H���dȐ��!(�;��/�uKM�ߎBB�.c��$2d����@��ڑ����䁇2d�~`Q�\r$4-!�0�dȐ�{�hj\���d�0).CȁdȐ��m�T�pU](�%ʐ����P\H�d��`2���HK��А@�O��m��#yky"2"�dt
����A���Y�C��w��]@:u����v<�N
��\�!C��
����r�B�C�2d�n��l��$2d�n�'�� �ѭPVQK�}��?����c=�|�{W�l����L5�G }�ѭ`����Bg3��V�q��Y����X2�T$C���3"�*R��2~�P+��P�ksOdȐ��6+(T�2d��J
���eȐ�,J�B!���wH�.C���dȐ�!��28d2�!C�L2d����@�2Ȑ!��Ǔ���<jht��+-����7l΢CGO�-,�"=���B
:U����O����taǞc$�g⇟w��	=�dȐ!2Ȑ!�C&2dp�d �Ga̘1Իwoɯ?p� ?~�?�8q"���K~�]�����z
d2�ѣ�h�"������I�/,<�\�ի���Iz��ɓ)<<��y��)P��	J>^�'2z
V�XA��Đ������h뎣v�>��3�����u;����SG��A���w����A���/���^$������4��/�?>�SB����Z5�g��*;QL�-m|�F���55�`�o:�����7�('���}:���J�C�uM�WPF�y51�a�;9�������O�FL�O�������SZj57��	���<44���&������08XG�}{��hb߷���}�}�f3g��Ɠ�Mˮ[/��^o톬V���|�T*%�����2��o��J?̑�/,���&����]T\I�U�'����JťUT^Q�t�ǎʠ��g�.(���S�Jo}Y��|h�@S3��z��'oC��?�>evT���?~I=^�	��2�-(P {�bTPu������7�Δ�!L��,��?v��7��3�3�6m9��B�HeM���8��z�	���D���f3z m�v�Z�4vL&�7���@�Fd��]�� �yu>	q�ԯ_ov��QS+��A�*�f�QQI-�P14���?�T�`6$�
�k((0�F��O;vgS����3aa���h�ٷ�8�^@��gPaq-��;�}�,�XCc�w),�e©fׄ�ߒ�פ�������5ٸ� <<.)k���q������i��m,�nY��9�Ե��n;s�976��51�?��s���9<���e�kl�!��i��cTǈb�о��U�q+�Heg��	aЀF@:��oadݛ�
%���8]��j
�a�ͿM�ܤ�T8��ģV�ǆ6=#�ꎈ�Pz�@:��j��T٬�c5
2��ɦ$2H
hF��2����;?�����q-7�N
w\2�Z�F���m�ẽ��+D0a�7���}��7��6��تh0bA����V��
e7l3a��oh�R��ma+y8b�R��jޞ��H���+�7��;�	dɕW��X�?9)��[fz��
DIY=��|����WB;�Ǝ�GE��:>.�d{-���`�E3���keBؾ�GEQpP �����]����+��B��wU�_7�������hf$`ݢ�ukll��n���E�UZ�����_Q�D����
��y0�}u/cd�+1��+bd̾s9�_�H�R]}.�B(�D�j�k�k2��
�c9�|?�mv��Ƞ0w;�V�QƐ�Y��5��=_3m�Cf��A�����dT��@��T��	5շ��M�d��Ng$pQ���1 �B�1��6WM?���V�KƐ+Y�g7��P�����Ƀ�4�j����Ps��i����+@��,lH��

���U
�&BM���r�ͩ��&�������h�pR%�iN�� 4l��J�_������s��#���U�O��|3߯b�ebj>����r���(�g�8������;�Ԝ\ ������UZ��ub���1�,�s�nМp=��-�]�|v��ta>X�[h��;�`���p�xƮIQq�zo��Z+�����WUW��g���o���7���m�|�ۅ�1�hry��*����un4H}MQ�"�J��iH�{MZ�^7>�D����!�)s}\�~��hd�t��1�̈j��Y����T����b�Ҷ��h9i�9�O�}�w�c6�ub��C�L�L�7|aQyǪv +���i��.a�iU��*"l�C�QFz������/g�@�ofDe�_T\�4�P��ú����c�`9�������k�������9\8A*�Ք�4��� �&�����'��';�����{�g��:j�H6�n�O]�&�m����mϾ�\�W0⩬��Ҳ��|/�?bX:)!��6p����0!T�,A��ye��?���k�66���ב�6���`��GQ���MB���6z�������Z�u�,~���4mt���e��I����w�6��� R�<��k��@\�]���}�^�-��fWM��K�����������C��o�ߩs��{�q��Xe���Z�rE�>Z�7G����p�刘5��|s��H�DTV����Zϴ;G��7lv��d㖃N�[�o�v�<!*��J~�g�9���Q��)TV��/�}�Ls�n��v��A�_��r	�b���]�()&��}��d" ��t�����L#U�(�p�s�ETZ��8͵:�hPX�je�a@�V��Sӌ\%��{�!�9QB�����~�	�v���^k����C%�
���
��V�a�/�X񺴔x��������Q�!�>�a6|�}O	���a2���z?���ܤoa�wE��$$Xǽ��t`�[�AA�<�V��rr�	d��(���Tl���jk<�ղ�&r�`Ƥ��n����u+��Ot5z���0�/<�7����S�{`�����i��c��3���N?��3�fґ�J�����abv�l��I�
5-J��""�@XŎ�c����j#J��E�U-J��2��?���-]�5wɂ��ODZl_��Oc�����`.c�G����܈����f.\�����0nU׶p�@�a3�A������ۦ���-۲x�m��Ljb�b��m�!���1���Le*q=��a�:R�Ç���QTTE0 *>� ���z
����B�f���#3��?8$�ƌ��r�������t���q&m�~��yT�}�6@˿�f���(�5�3R�Q�xv�6o�b�����U��n�n�2�Ե��v���y�A~��uӛ��`,;���u�)�
u�`������ɬ��NݢG��.��u�X
��,ر���clӳ{��t�ޝϦCy���������������Z�T`e��O���W��;V��m�sϬ���oY��W�԰x�H!2@�s�M���\p"v�`�D���ǵc~|c����޲g��a�⯆���-v�?$�g��Ѥ�G�����>��~�w���hŒ9�V�مt�_R����8Xm[Z��~m�m�p��Mj4	T[�n�j�ǽ���)�����r=�	5[�kڝ\�*��u4!������\`�B�G
�
��!�zz}[�m�;9�D=w�a�8MH��=�������hB�nU����#�c�ʏ�%Br�(@X�����]46:z<��p��*��b:u�Bگ�
(�-���56:\�z\�H*�^����VY��Q�/�[g0h� ���,��cB�Ӊ���#<�p��u�;wl2w�J4�{/�H�Ξȅ�ݟw����径�|��>��s�Hf�At����*k~<����e�u�,me��yK�[3>��9�C;B�)�R#,�Q����^v$+>|����s\��߶��H�0Sv�{�-1*�>z�2�,t���A�f~��k�z�]�?_:��d��}�c��UKk�r[�ө�Z��Lk�Ÿ�	'4 �F�Y��롞Cx5j�������L  ��6j a

�d A���p�E2M� ���؟�ƅ|$��!�oBH/��ǹ�{�M�����(��P���@ݩ����*v@��~蘈2�����uk3�_7�z=�n&��ҭ��������ƍ�7)X�jUL�2�(�}�n�y�[��'���'�^�a;=����z�a��܋�?�L��#�ӭO��H��Ϋ*,?��_kK�X��U�Y�[�'���n��V�� '2@҂#�̭6-uw�ʺ�'���92P��<✁)�+*�.|�U*�m�Ε�L3���zU�lm\4$&��5�=���-oϤ�+(�Ysr�i@�d�����#3��}JaYyuG������U�L;�'o�h��b�y�l���f(��GK����=@�kTd{� �kx�����D����V'ceu��6��S(�p.7���XSSK��㹴f/�����]����'�;| � ���[~iG����VPX�|ݘ�����nY�2�\7k�`W����/x�W�� �B��մ��)'/̄E�~C?�8J�F�����9�Ai��y�+�q���V�9�g��>|^�V�2wd��BG��Iؾ��jw��k��zr�I�4��Ŏ���T6���5���î����~i	M.��%Uv<+�y��mp��{�ٰ��ݵ׹KVd"�>1:��7Gd��/��s������_P�7Gxe�`׭��׭;�SH����u8�#�� ��_����wg�M
t�}�"��#b9,��Q6�Ƞ��,pAA1���36���˳�}風 ���t%��L'��CSh�|�־:Y�߃S�O���u�0~�x>|8��ـY�nݺ��eO@D�oZ2�誘9���H���|�7ҍ��-�,"���.��+'Q��V�d�/:�AU��"2�/���F�ٮ>P�fY�)�n�<�}͞c��X1���ژ��l�t�rse*����.?���iG��p��Zx�~����O�3�<C�ׯ��z�ZWV5r��(�=�ٔ��� ��F&�%�Jٌ�h/�w��_���K��D����i׵�ω
�\;�ګ��̗��_x�7�/��=7��ec�8��q
�=�A3�Y�-���5oű������ǿv8���H˿�H����$����ԩSyh�R� Y�������ʡYx"[�K�&�I��U�MTZ���H�"�~,�I����mX��3N�[�?����Q�����(=�@�v����0�NE�i���^xcM���=���9���1$�p�V���	����&f�����Kg����e�<��Iff&y�AHp%�������{���V<yǥ.�C���;�y��U1-;�NIi�R$h��3�IZ�`Em��ʢ܀���1!��5���,qN1M:B���^fz�"vcMS�éӞ��P�
m�59�ӑMx���(%>�����[EY�e4}L&Ϳ|"]���$��(�5���ѣG��>d}�8X�`��k�X�x���A/9��cj�w��#.B'���m��@�Rf{d�U|��AA{+����Ҋ���м���������Z�=2���x�۪	L�No.��^�z-��bZ��8#q"b����(x[U%�G�?��|�R�>�fn	��u�u*Z����)�-�mL�>�
-"t�t�/W�7L�f�7zE��/�tĤ!i\#���7x�6�������x~B/ϸ���w&�F���X�|�b$�g`Pfo�����+v)�Ef��i�[���4����	�����Ri��@���cTӢ�ky�#O����#N$��zj�6%�5'�ei@*�?ڡɐ�ըmj�م��phP�d���j�>z*�+x�PI��{4�0����it��b�=���
��4���5�W�O|��G"hj1R��� ˮ���;ɐ!H���STxPGj����[��̄��&WM���]�j��q� ^Sܠ�-�j�^�ٙ/��_}B�6�� ��t
ֶ��9��&����8��'�/'m�9�	Sx��'?�ͮ9�/N�^G�h�������-崵)�f��(j�!��;!�d�p�}�*he^��eFCF�_H��%:�.;��>:I$�ź�Q����Z��QB���u��	��iO��l�u�~Us�E��Ha��)�������R

����T���ې�
�Xb������"�����}�[�J��w��#��l/�����&�(7���v�02:��,���J(-�T�5/+��0|w^�X�a�xNWp	uXH��.T?�PA]���N��KM5ر/�ƹR�V���RJ��"8Z�Ȉ�~a�V�Ul`dpj_NI�=�R�E40i	�� %�Z{eG�t�8�(��B��#�X���Y�e��6&���A�ݾ�Ӕ�uD��nE����#��B��7����F8��HG�4��}MP��HJ:VI�O��=��44�����sz�_�(��\D����d�PFp#MM2d�Z��3���ݗO%m���ӌAZ��'����9�vOe�DSy���A2�44�L�-h!��o6�&�R��J5��'��-ni���D��L�a����whQ��z�a0�7#��			G!!!�������Д��jkk����jjn������ �鼠���6���hΤD�u��>,83d,�0&��Q
cr�SL�OT�br�U�$���J� �.N3�y)F����D�!����L#m���Ϲ*Iܓ��v ����uj�5k��ĸ}͇~ȅ�3@�W���y}KmL���ί������:���:��ޕlV#��7;e	C6���<K�Ѡ��9j�R�v;��-D
t��
�\�	���f��1fzk��k�X#B����K�yoW8QPIUU�� �m�2}�t���Zӣ������KG���T�(11�����0��a) r������b�~��#�d���B�%��v�56�7m=R �m�/��ɴ��Y@�H�2� )38T+������4.k�d�>�ϣ|��7H��=c�h�� �HR1�Q���/}%�W��=:xr��#��t3Y�_���^p�I[�n���_~��7�=����@:��s�o߾t�b:t(ߠ%���pR�66��7��d��IB����IM�Ex����[?P���ht�z򎙔�M�,|�W/JAr�@w�4���� ���)Ы��$�P	*��ý'+���f��w���`�~�Ŵ�`.���Mǘp�s_���@5�x`/o>���H
0D%�]`����ԓ0l�0***��;3lw+�v�� PF���~��Z�%�ps��Ȁ��!;;��9���j����V��q��(���}J��m:���;i����ϻ�3�����t�ޗLo�>��4>Z��(0?��cΡuQ2��0=R��Z���YQ�S	�Ia�L���ӏ�(c����:!2��S��p-ń�����ｒw?��k�O~�O��"�L�0~0�Ե0ս�g��}��ܝ�@{o�d0mڴ�jkUU/H����'"�B�z��f�!�֪�ç 4������l�/xZ��5��o�N$�j0@�����M`���`.I���'h���A��">f��'1aV���m����[�K�E�&
s��Xڤh��+w�,��`��j�%S'2U�m)R9�$%W����UG��'~�����w/�Y���8���_�N\
���MO|D�.�C=|�}�c����X���m����qM�x���Fw�Knr[!�`xr�!�e������'�����y�vƌ.������;Ʒ�j�͵9��ܪɠU��k3h�ĉ��@
�@��X*�l�2����I�R��M-����7:�K̂I���[8Ė"�g+B#��cK;8g��~�c[��[�<�j�3���L��z �I�	s>��je��J��ʕvg�򥥸{�>�����FXRl��͎��in�de}�H�_0��:���O�A�-��w�mi3rA
�G����]�M�:_���`ҤI|����+ݗ�B������� <�~�,l�9`�v2����ߧ���|�s�9�����!v�t����c�������T��}Ĉ����I��^#O�p��iD06#����R��'1����{�z��t���|�:zyBf�E�O��D�ۊ��_����?q�#��*��;}b�����ؙ�NW,�@�R,q$[T�(ocd��v���-u����>]G�̹�n�d��s�{�p5
U����������Dn�_��=��C=������W^Od��Izz��~�R9 ����� 2�|���PXT�M�W�u4�P�?lXZ"�|�&ڟ[F3��e��?����ү�|x�����o�h¢��C������D��"�5�޳�/V�>�୨@�m�c��
vU�Nd&2Q�Ũ�o+K>pw�o<����O�7��2�j���+�~�+���P�&+��W5J~�]{��,2h�[+8� m�S���5�B�8]D���RRR�& 2�ZIg�%���m��D��)�<@H���������ێ��^��u4�q�0k��QY�룧�'�؀���ϟ�#��-��^�0x�@TX���J/��w�C'�'�߬����l6w�����qz B��ʒ<��߰�����:���^�����zF�օV�)
�Yώ�"nf�ͼM��C�}���N�=iG�t"��� $6�.����/]}�m>8&X������ޱ��_���	����Ә�ω�o�]ST��}�S�t�{�_|��c���s���N��R b�K�AfzͻAZ�JY����Q��W�V}J<Ex������3����Xvo{$&K1�����K��]^L&�z����<'2(j/��-<�� +C��"um��/j�V�D�?x=g�e���%לO������է�f�6l{og��C�{��ZC�N�����X�
%����lN�YF�"��-&"d0�w'����5��^w�0�c ������;?I�V,"K�ZR\k|o�Ub�vѢ�ޑ��#!��� �Sz��k�c�}np���u-Sv��Z�ڱt))��|�m�x�Rv�j	-��[���ps ��CN�V,����T��=\͓!���O��b�L@΀���/��D%'�>��&�ٹD���{$�p��g�Dj|��J�E�>z�%���X�0"-̼'.����%G����V��?v6E�'�'�	h���_�f�N#��44ed�Y4�l}���M��+���P)�`V2���w���r�|t$Oq�փe��,��B �T�U�B)4DZ"KO���I��Ƶkג��g�'��������E����n�������&� r���Pp~�ҷ[%�jT��b5ML���!�89Ÿ8���R�W�5��@�bhJ�y�XB |�$f �*Q󤄤PgBHt�!���w'^Ԩ�������׾�����ky��g�7�SmoN%��B�m���q_v�,=լr[��VF��|s�i� J�w��E���\��=�7nt��y�x�Ф���g�m�ځ0j�׸B����6����u�ET�=T�cs_���pd��D�r�K4ۮ�t�m�P�f'�J+���}ZZ8�ͩ���������,���|�3z}�54~@�o�:�?QZMSz��1�zSsK�Z�v�8k'���������� b��������0l��цT�s�rb�k�9�����щاO�t��P^-#�n�h��'��.�!�Eu�z�=�5��e�=N�=v�t�a���J5��g�
&�w�2x����W�⋴˥-�_ݭ�ۆx)�TԲ�}l�C�����е�y�&JqzN�D����$�4��D$������ 1� kʱ١l�-��PJZ2��09l���lU�j�X�{����s�a���"��k�g`昼�_Kb �����.#��%� �˷��P1��[�:���l���+�\$5���
	��Dk����%*�(1�wϱ��Y{III<�G,�jvii)'	�њ���$� 5(7ޱc�L���Z�F�H�q$�H��!��``�pҕ�R+��+�3�c��N�L[�'�P�H��~?G��T��+2�.�
��X�u�Z�L���h�C�?:��_s-4"�̛�D��;h�CT��T�h#�2��	ѩ�P��uc�c���SCk��I�6
�TU]?R�uQNg�TYT�!��	��!dؐ8��~�5�a@Ga�Ɠ����X���jCG���d´@�-�=AdR��]H�eV���AT.DF��N������ �9���Yz*6ǒ����Ѻ�wp2o��Qf�ԡѐ@��Sm������s�����O`�~-��QI	1�;M�H�#o25��8��
��9���B>(�pA�^�n>��|>'�� ��h�MU���
�P#|�^z)OK>�����DӃ}p�4���|����iQ��Å�Q�g�?8^��O<�zDwd�DAS���O!�y�; �pgm���:���v� ���&!��ĉ^U�����yM�-`.\��\C������ٚ� ��Q􀼵A�˚�%�A.�o���+V��+�Y@K���͝>�l�0�=�����Ǟ={xYsw
�:sg��puYm$3����Ǟ����@�-��2��jZ����N<8��o�Uw�!C��Uv�Ν>�ߔ)S:��d�6?���+��R�^@�1c�pEw5-��������{ ������&}��l'1`���݄m��:��0�3@X��m�Ɖ�u��j:އ$$��+�5SP�m�@$�4� x*a����'Ԁx[�|6�k3!@��$i���X��n�n�!%'�Pz�dv�Zxb�tE��>���>�� ��Q���F�A����G�V���"������駟�l��O���EʀG@�={6�X� :�5�V(�u;:�Ԍ��onRR湕[W	��CT���+d�"�F`r��^&�`���]�2�NI��Դ�DEg��~���zӑc�m���y�䢒*:��
>r�H������e�IjQ�cA�����￧�3g:���}5`
�\�ży�$7@0;� �P8,��d��ɱ��&P��NE2zSiy5�鯄n���6Ѱ8S`$�Q���C���2�wfZ���l�� �ob@�徑������)����N�f�6����]0qI;b~� }Eo�dx���^������ ��Vu��-�ܭ�FR�ā�����!LA8�Uj�C����J �3�ݰ@#!0���&�J��S����\[p�d�����J&]!&�Bc���Cw�zGH�D�(�Uf��|Z�V�'�d2SCc�"��`���@ڲ=�N'pSX�l� ��ꫯ��^�x2����� 9�9t��
d�A3�kgg�(�=@Rf�8�4!�"9�$U�V��E�TS[��Aj|$�r�h��k�"��	\�"=��Fo��RA�����fo�����s���F-��F������a��X�}����A��1i)<8���z��������"؏@G���1�� r	ۗ`��b�7�~�,�ݏ,E8!܎@]��}8*�#�2��c�`f�	3r�h�^b-�7m��#����<[�g�!*҇�x�d�u�Xz���u�LI5yEV��p�H-ߦu�� ����7���� ��M*j�p��F��D���o�)#iP�xz�ˍ�����t1�|��=����Wt]�Ql� 
�7g���`6|��v����?P��4 =x ��>���#sp�رNQ_jC�~���!��'���W�}K5��Њ��Q!��XWH
hf�#d(#���&Ҙ!z��EK��<\�:Xьh���^(,m�v ������e��,/4�\�+��4xw��y�'��)�[��a6���q�ec)4�w?Ŋ����3���t�G�c���h�Q'�k���7�����H8>�o*����A	�9.5 C�|g+0$eS�}E^-�f���Wtm~�n���\ʈ@�H�&�p�R����^���irB��0=��Tc�Z�9j�Nd�s��9VhdD�6G��/���6�aȿ7w�?��l|�qd��$3�����qE�3���ĎB�w��ѫS=?b*Z�Nb&ls1�A����BX]� �㪚�/��8�j8����rX����T����gH܂�yۏ1<,�F�H'�q��6��}�~��׽\�����n�}��yC��O��CR PF��lַ)��r���56�!�O���J0;5D�$�0~=Bdv®�oDЁ��z���[0mD��J���΄nI���v�x1�6��[�_K+�����6}HJ'DP�,u8eWC,1�!]�r����r�Mx3(��/��t��z�)��Ld��� Z��[��"C��r2ؘ���\B��El`�Y�;זb�R"��+�}�/�ob�H���m&h�yNd�Lp��(�;Q-�c�t쾂�5�[�qɍ���k��չ�ڞ%\[p5����f]F�M�X��u���j�o��#������~)��^㮯��{��Q�0��nKr��D���s�[���}�T�@�6�:��Fa��=�s��WM\��G#�E�~Co.��wF�%�Dc�b�8��~e���Ed�c��Wլx�o$=k�MQ�٢oۄȉ�|�F���ͧ���{���e�!�n��:Q	S�0�>H$'����m�%ǔH9�ľX.]~�}`AI-�p(��B��gz��|�{�xI�/���C�p�a%w��h" H�3G\}�'�6�P(����?"R���L�31�@�t�ԩNu������/n2S���g9L!���DK�m��SD�㿶��rM���a*7=��`��\qϳ��UL6��PGK���Di�?��G�x5�d`09/�*R�{ۃ���z�e>�ҥK��*��I\��D�g���pV�v+��%4I�ԔB3��L�N�B�7u�{�RhvC�(��1�)�bف���!81��ED����Ҙq��.aM�.@ �D��D)d��bGX��1�B���bZ�ѣG}n���[͈��7A���#9t�Sћ��ZFI��{{��(*��~�)����6)Z,�_�<�`M4 t:��2�$�u"U��dJi}�=���,l��S�HgG'j<���/��G������0y8�������GA��L��М��z��=ݨ7���F���;�ڜ��;���#.��Q ���G;{�!�]�+ B����	ռ+�t�"¯��@�E��W4��/�������F��7�OMr��q�n�pO��{�׭�˒�P'!S�z`�/�=�2+�	�|��umF��թxN�������@ɟ}y�+�q�}/��Ñ��'��9�&��p��t�1&���}��>N�࿷N���x}�%�m�8�q����t�a!�&J��_gd1�����#G2 \�(�U"1	���q\}��j�!�Ѡ���ɫ���.$`!��@R���A��
"U��I�̌����z��&�@F��z�"���#�_��7~t� �s�t>����w��p�VI��AN������kSĦ��t��3�3��Kr����tGBAq�m�b�^�Ԑ�����}��ӟ[�߸h����������2{�Z))�H�m_	1��P�����T��L�ӍC���{�/K�逡=�J�tcFF�mҼ�t�~� ���������OS���>t�-H��d ��5+@ܰ����|�:PCK���Z��� 1��BgM���0�2>��*�CF��Y��("�2����B���RZ��@�$��&�9Q,�<�#����=�
15Q:[�5'-T��;����~z��}��s/Z4,��N�(w^�D���'4��t��0!()������ע7Rm����B,�bI����q͘��ͩ�4�o[U����ȷ\Cյ��4H�c7����
T�9��j��_͝b�Aw��EJp:��)���v�1�`k.������>)xk/F�*m�����y���Ӹ6G����D��!O���d�%>�_�C�&���&*�j���`
���GS�h��bZ]sz�� ��s������6'��P����&�B DGEM�7J$�b�Bl*PӤ>��:�i	X~����\���ﲮ.��[�9bD?����y�;DG���N�����G���ӹP���ؽk֬�q�y牾�-� S�K�&�ʛ!җ��#� ?�(��g�| �h�s�~6�� 
�S8"�j\�����:��^	�ӷ��P��bB���&���A���l�K�.�|[����RRJ�����w��Ip�\��l����r�>����'O8�̌���'�Ԟ �ԝ�\�*Ts[�u-�X��l��ۏ;
;�[k)2�z�׮Th��(����D�~b�: _:!�so���q~�i�V�9|�����v "�"h�ڝ�iI�3X|��._��ZJ� � ���k�H��ZЯyj>�D.� �=o��r�dl/鄰�DM�Q{����}'hȟ��^UW���d���?���{o�&�z��fE�N��j[��Ŋ�
���=bD�����~��7�d�`)�[|
Q�d��>u�x1=��>��ӏ��s�t��ǧ;�oĀ�I��a�ڳ����QA �o��[�����/�h��YZ�[n�KӍNc�mQҤ��؇��-����ik����@��ɱ
z��
��p���Yg�\�:x�,�
�@���U4�
��	m	N���L���վ�C�@#�
�s���Z-�tN����599���#���>t�$�8�HU %[h@���^Df!�u�
��Jt���ĆN#�FM��TXT�e���� ��bN�� D��$JVXD�	�P��p*�� W�]D���B��ݥSRj�x�Ǜ����T��?������jގ0=�L:��ĝ��z%f���t:LU:S#Լ�葙�_X˛��MMd�e��u]�nشP���NE��"~�c�� )@"|	جݘ�P1�qhͥ@D+?B��R��3�a����0JH���U���v�m��9+�+ R@[�����f��b-�p/Y���5��+�  !l߾��n��(B�3�Ǚ,�poˉ�#p�Զ�)� ��r�y��ǑH@ Oc�㘨`�w��|���>�0#�'�|���#��c%>��L�����KM�6
�i���ID �82 v�ʦ��R!�R���o蜳�����K��鈝�ݚ�QS�D��E���Ζ�6ڹ;�zz$����]�B�-����� �g`O�DJ�j��S� |1 ���n�S[���A���t�����f�u��.��� @)1ڭ�Z��*�$!oS��
��a4z��m�*ML�3����E�)��(�!��e��3٬VQ�DѐDHl@G�~�NBp���)���^L�՘v��N�@ܼ�L>��[����D$d]"Ԉ�BW�g	�t�l����VP��	��dqD����3�v(���_��Y��~�vKha��-��qO-8�~��?�����c�s)e8 B��fOs�@�F�}��~� ��!�I��a���P�32�LCi|~DKۋ]gB�$p�ܡ�]m��)&�
��}ZɄ0ip*=���h��yZ��BwN��G��[�^IM-�*����4�}nJ�x%�^�ƎQCMl�����)��ʐT&����Z��XmK�Q�4a��)���vw-��:��B�����b���������Ԥ�%ǄSnY���GTRӞ협C��u.My�5���F��v��V������A
�jhM��ػ$����0����;.�%B1a�����+Υ�f��7�A�K�(0@K��:�V,�C���}^����T�zH��j�h��^-���n�Fj//]�~��U9t�h��d8-�l�0*�P����n#c����J�O R�-YW���ՔeHm���h[y�;9ȉ>�\A���5	V�����y!�_����l"}�7Ҝ�>��»xEJ"h��F��b:3)*���ܙ�D�iǓ݌o�mQ��FES�V��	��89�H�˼OS�>&�w;���V���Vz�Kم��Z�p���2ߔ���Lv+����oi�	�\�J��[��p"j`�A`�34ۊLd"=u���o�}
P~�q4�����BK�8���XQR�����})1*��?�&.��s9X	�[�J4Q�Ġ��fe��,�Fh)4$@pr�Aپ"��K������lUW��pY�Ұ�B��g�yɺ���#�l��o��_��H+�{�़���&F�M�m�X��&P]C#EE���[��\>�vV�5z��V<�vH�EA ���!w!5��j�Uە]���k��a<���@w#+	ئ[M=�Qm����؀���W����Z��'[���_�W^�I�J�~�Q�y�H����۱UՑj͜o^X����t��oE��[�ړ���MN�Nd�	�c�Uq�g_�g�����"(�?��[X�Z��΍���:����n���x�m�$��şv�Ը�v�6z�Lz��/�I
l�\�>)!V��/@�k�"�hTbz2�����r�A�1�b67��vժU��M�4It�o���KB�ꪫ�2Dűi�mR���2Y�M��F�hvn"��"�� 96���J]�Z�<�����	�z JE�p�h��je嗵���_Xֱj�[�Դ���/�mB��;&�v'9"���"�f���r�s�D`�;O.-���������)*ƭ����,I&1�-��;{"'�;����/K�Wmt;tU-隴*�ٷ�6<��7հ߶]�U),tyB��O���nt��ЪZ����Q���`K6�bl˞]���Y����AjrM,ȥ��S�Wi�ht�����������Lc*�8!l:����*�h�|�ߖ�: �!#�y�6�K��Jq��U�?xj�Q�޷vh�e����a���Ap"�� �ĜŃ:��jܿ�h�# �����ܓ�����Ͷ��M~ܙM����-p���5��O�[|M�̡1�B):�y� L��'��`N5�
�?)�b�C��D�2��!���w�ь3\>֭[�_Uz�̙�uTix���A�dW�2a	��`�L�/�G���l�)��a���	 �(tN�u8v��˫'&Ш�b*�j��pH�ͱ�dL"dZѦ#�lv��qxϋ_҃�^�Ԝ�p#��gM��*��\�"�Yڨԯy�Y�����z�Ȟ�]0F��Ƨ�D:�{�ͤ|����,]���ԓCM��CQ'!���r/�`b��V�0*-��8tU�O�֌:�4@>�q!P�!hh��
־V�
��P��y�aB@�0E�9 �cH�H�f� ��o�����^y啼����s�yC�NDf�m_��;2�.HcBZ����I��ʆ
��"���~}�z�{I�#*�f��		4����ԸWNE�DT��ܽp�֗�&�k�� u���6I�������QJ�s� ڢ���/�����ۭu�Ȯ���� �	��'X�"��-�����ݤf<��7�x��)�r��<��9���\@�V2���:>!5�;�	�Ʋc�(f(8b��|����%u�ҋ�f�V��	O��564+'S��"�h�0D�����xz+��TT끴��b�+�=�zE��Ǐ�@mL���W��4j�3S��\t-�}�c��أ�����7��:�Ԡ v��l�j��FL���õ	���S�@4���u0C`VX#8��tE���V2��uw�V��+"�EU���?���F-3Q����|�ȍ���>]�$���e&�g������ڌ��J�t�`As�=|������X����n{'2��th�=�F�2NoX���/�}�%��̻��A����-Za�g2?�w�L~�U����:==v�t�gP.Ҥ$�h	Y��\�B�:����)���/� :&C�@r�sW����<A�D-�w@��њCP����:����C����@������p��AO������I֑Nd����^�'.�f��:��\Ǝ��{ǆ���� p�REWf:�ЌK6?i�w���_x�i��-x�_�٩ә@�p"P��5MI��� �[OIi{1�7T��ʭAJ��������)��C`g����O�7V5��իO�T��>,4$���˄D�V�
��/�Ӊ�}���qh)2�8b@^T|lP�!\�<5;���� B����|X��^�o��v��� h7R'!� ��O��㻠#44$_�v'�KK��^�d`����\�7K�3�v�]h��)��B�L��9��1A�zJӶ�~�ܦZ֦0U(�ǆZ��e(v;�(����K���I6�h[ g`T��\�����C�QA��I���O��A'���j��>1��kj��(��}���\@�	`�0G�m�Ā�^�HD�V{��o"Ti�d�_1 l	[����(���V pp.8WhV����y�X���֓�^�Qt,��;�G��O6u}Dt GA�����	I��E_���L[?P!� ���G��f"z���5N�=CTL"����atD6�N@}C+EE��62� C�0��6r ��ꫯv�Gwb�8��H����ʻ"tFFF�G`u��f���y�|P=�ע�
��
���iF��Ʌw=�s�%�"� ��r8ym������L�$�O��$�Rr�C{�/�h�F�������\ERq ���ȥ`�xVZ��H��8�v�Ɠ=����m���ڽ��N�!@��x�D���p��T�����~Ǳg��AF14k��>��c�4h�T`|����0s.��B���;�I���2�3��[|�40)D�z�����F����o���*F)��iD�zyG�l�g������6`S���[�t� ��!���ؕ�4t�J: �J�h����}��هb��(�p.��W�v3�nl��#�� W ��l��]~�NBk��z ڂ�a#�1g�O[���.����@�T@dR�����Z�Z�����o�1��hv>���h���H������~�O�0EA3ҍ�|��`�����Rp�)A�ߤ�I}�4*�B�"S�P���TM
UN�3L��w ��
�6��Q��P�ZC��W�`Rkmރh lmO���|�M ���@(��V�'Z�ä8:B]���=�CrEe�i���@�5pTM0S�Â-�Ƕ��|z��$5@��/���W<E���	E��g��!��K*��mώ/a�o�``5v�?��y��aBh� ��J���[�X�m�6��@ ,���
B|pvR�	=	!�:�,-�R�A�t&����,Ǡ� �˧N�>�}���
��#���ۼ3N7n�fb�z .��[���[;u����jk;N:x�Zt%\H�E�	�D�!ja+z"�'B�P��4gD'@��FRp:4L��i)�4���}~?z ~��=m���R����葭��`�Ϟ=����K���"����+02a�  8B�����]4�߆U����B��Щ�,QKڶm�h)2H�S�1B�� zҝ˙O�dp�DOA:-� �����jl5Q�^aH��o���
m���?�9s�����f��s!x�@B���D$>&
��x�Ay[l�. WMTϔf ��F*�j��H%Ǉ�|]um�-�;;�#���4����n�_��촭�H�nj�|s��_S`��SJiDF�(B�:M�2���l�z���7rM�j"௵F �M��u;BҒ���tu+�v�y
ؤt7�.N�w���) 9�ʣ9�:W�n�_F�T��Y����]�#� ht��p�K����yo5#�SM*�����	4(����H<�696 �>)5j`��{˚ � l�������q���}��<���JP݉p���u:QXVGk��2"8�o{3�>��4�f���ӷ���O&��Ҁ�Ű3�6ST�@�����T�x��LG�0�m����S=�����JTZY������Y�HF��R*� �B
�\�]h�Lf�`�DJ� ��i��;�_˫h��˫��p��*�d�3�v?)��;��fmѐw�hh�ΪT��
%O8��d��4�����m&���5�H��cBk���*�!G#�O��,,�>F�i�\����Q���`e~��:�����GR� 	8�`f�9�c�#���uw��mD ��J�hRs���FKJ�4�Z����� :X<Z�9zfjo:>���eF>���+�6��f�'Z���j��LܒAL��nip9���@L�'�1sbxk_�W!S�G�'�~q��hD:�G�ж#�t��}y'0-���*�yS����6�9يI�y��g�� Ƨ���W�
o�Q8�ܑ2���_~9�q���a���Px�����U�>m5�t��BG�C}J)�t�^�U����Z@��H�]H������K���Yy<+�!i�ly�����-2��4o��-Ȟe� ��{�;�u�X�$�3��X�SV�'�8��J�n�I6p�����i��|�h���i����@���v_���^DCҝ��E�ђ1���h15T�+Ш��'�U�}�#� ���1� a�1�[XUsx�Q�`MU���_��; � 
��cW�����Ci��*hPQ<[�%�c�w~4me��]hG��s�pz����'J��ޚE�N˟k5����Wr������EZ�b@���a�Wv�I��%��7��@F���3��8�7e�ӑ�J��9��\��A�톩��{i���ꂫ��%�Ѹ/pbp���:�IG��0{|0��O��C�!��ʰ��~O�F���u9* �8��L:��@�ʳ���f��t�p�S�@��=ZA9"IG��9|�� =��&ޱD�� �~�����rz��k��E/RU��ķ`�	�2�{"�Dri��g-:B�0�oCu��Tؤ�i0�rtKJr�06*��5���;��s�"Z����;���?LNG�*ُ��~��;��.ګ�]E���dp&���Z5hVK�7N1hR�j�
Y�����.ߥ3�=���܀�ԛ4���C#x���2]��m=��7�(�ů�Ї��"C�$�J�C��OQ�R_�L[,EU�F�!c��D��6�"D���d�j���R��'"&e�\����1~@z�j��X�$��_�j�D ����t��}�%\#��G�V���a��;�B�jП��!`��`�+�G�S�M�:�B��(e�֭��	8>2&񙨥���UY:���X� ���Ǆ��h�L����~\��|Ei���)_��`._��&�H�J�	��e�6����巒Mc�k-JJ�0�L���b�*ŀ�/�k�st%�9߄G��e��"F�ʥvO����h�xރKK����+�'�w����ت�������贜Y�=��[�&����hD[X�d!C����p`���F�� �ZCs����p็��HAFT 1�iӦ�<O@ |RW��<���� ��ч�NP�p#����J�e���7�}~�&y�F8�/�m�M|17�wqU=���V�\`���<��&ϦـhL����Ռnqܿ�g��}�!ZmYlم�eXuDcg�;�Ar�EtXDv��~zi�K���ۻ�(���nO�J�KG����YPE==OAP��=�;==P�D�+("���{	�$��޳�?ϗL2�;�;�i��l�����|o}޼J��Jۅ��8	�UI��.���g�󝃻�i3 d�zw9U������Њ�z]J�n���	'N���$bW���j�(��*Q��ߑ�s7�	��;^�@9Ԍ�����@A$�ݱ��zp�H3���@k�޽���\KnD@�/%���
�zLI˖�NA��%����g.Ӳ-uV��w���b�y+��
�:���ʍd=�r��׬|gqq���-��3Oޏ�� ��(ȯ;�A��,7ȗ��
t����;���9�Y���lV���\�0c�Z�i�)�i�u2-GT5Y��51���,!_� �/���?M�~��@B�1 X����&� tJI����0
���9���6&'�K���Z���[6��n��2IH$�TAJ�8��Ӊ�3���L}{����H
Vm?N���ذ !>�x�Vn;Fgӥ�uA>��Zv�����9.�b%����:���ҹ!��Hj�Ll���t"�Ƚ���*�U���Qi���RB�F��b����.2���￳8��bӉ� v[ȟ=��C��E�}��� ��ܰ�q�hRr�F�5��:W������o
�".6�2�K�����:���(�y�a��8܏�N*D�%���l@����ϳC��D%�St7g��r����zf0�<�Db�0k�"na?��rJ� y^V^�-�0*(,g;��M�����b��s��3��Ft�R˘��D ߨATwY|/؍�7E v|�v����X>��ϡ�5����iR|��m7nl��r� "#����ŵp�J%�q���OO`2�㺩��Dd�OT�5d��iA{�Y�4SE����s�M�\�ddc�&�­���=9��Z*&���À��6�X!|4j��~�~���W�#'��"#B�cR�ѓ�.�Na��\<o���_�r%����+?�*�`u`�oڴ����p����Pi�˭Ad�v��j��(�FB�R�0�+�����,<�<!  �4���+y����
+�x���K��hF�r.�[�m�-������Ƴ�/.r9e[KRt�Q.�Kt��k~x�b��/��3��*7d��F��5?�5������m���tN�~?j�uwc�Ƥ0sG�c��*�PB&�ud����wь��?�`u�~>n� H>�ʑY*5`ׅ�Jp!��
ؙl����s�nA�	
Y��RՉ��y" P��]��-�RvZ9��Ŧ s1�F�M`y@��1]Ml��\Wq���"x��(#�q�~w�VVg��N�X�}�ѠX�X��3-���f�?<kVT\��P��šL�C��`s������k�\P|���v����91^�?,2�*�ݲ5ճa+y�z}}4�+u�-*+ff�8��c����j�*.b,N��G� ��Q7o�,�:�k�
��MX P4BsjpΨO@�f�Tu�"��q4i�U�U"Ĉ#�e�O������y�x�Ը�n���s��+j�`kqiTV�1��T�7�?�]��fUP����=1�j@��1�f%4-�Ct��Rш%%;��Q�m�?��xz��O+Vҡ̦�J|�ٱͪ���!!x�����:�.�+ 0_ʌv[WB � ��kޚ�I
Y,4��.@ReȚ�@P��+ĻN���<��A `�g�A�N��	�_/��o�Y�Ȏ[�A�m��c캬��FBQ2��,=����%�K��Y��^/������w�<�U���.�S��{Ā;4|t�Bc���.�� �e2�i9���2Hρx�Z?�Ij6��� ���of�#��l� q���;&l��˅�Fj̣)`��fw/x���^�e����[[O��;H
H&2�='n9��`�䠖�cd��R�_��ώh�P/�L;|�f�E[y ���dxeY��܉NU�T^a��� jH��߾}���]�`a�U@��G�Z# "�� ���d)9w�՘��� V�̄b ��R�ׯo���`�D �Z��W�f���� ������ ���������_y�8�JNq{m�qn�}�+\,Tr����'����%}yL+ڱ�<����WGc�4(��r�����*Z^��ET���^��><G1��hJ_E�ٺC�aO6�)k���"���QI�[���D̥��`*��R�T� ��@ ʎ��]&6���=�%��`a��.@*3-	��>ˀ�'F����J���,A��y��>8r6�V�FQ%E���tG��ӱ��̥<Z~!�J�mD����\��p*WI���ĎF��:u�Sޜ��^���^uJK[R,Ի��:����
Z)˹7)�T��KG���W�|Zp����p.�m{?+w����}ʣ�ℂ^����Q}��ȕ��*�2�.�����>�FX�Rۡ��#�����+A�U�Є��]M����Ea\ �[�,�A^H����ρ��-�v�<%�����a��`MV�ˠ��u�j0f�� �����Ň�,��+�L�,���Wme5x<9OEG�Tl���d#��K�]��W,�TRV@Au������f��`��ͤ��P$��?g@`����E S�?\w)2��"�𥑳��+V8ݵ���A����7�?��A0MX'Ȣ�����e��)b�Ca	"0 z2�9�W|?�|����I/����U��n�Ƞ%4��Y X�[}q��l/�D��N��G)�+��F�-�nD�=�v,B᱐NDA�+ �����X�T#��T��Hp,(^��θE�Uhj ���	�����l��'`��dK�O�*�����>N�C�%�|�-C�G�"��~i��Cіc���j��tҤSx����R�]~>�r0Y��p�f;�+sZ x�>�&1L\wd k��ֱ�k� A��c����$i����K-b�/���?���|�\�(^!.��G�@\@Hx �'��BfEH >��dн]8�])�kݮ�Cz�d�7�.>����2��%�E�A+e�.�1};�'���˴9UC�fu,���4�>v)��X��&����;�5��E��w���Fx/� !�vQO�ƱH�^�);��L`��]��`] �/�p`����?Lz�x�i	AY�@PhdOp�x2�g�Wl��'@c�3��h��)R]A�w�R�]w*��'kh��:]FED�2Z<��B�����:���n�o���!��O1����w�ۏE���/9�Q�/Ʀ;��D���G ҕ�����}��Q׀,�x��� ��Lj�Y���`�`�<y�L��D7'�d]��,�n�CH�-�	���ymt?�σvƽC�k���32��5`fB��X�
!�W`�Ctf*vD���� ��D�y1R �-���`! P(�S`����}��
���b�q�_�% x��9r�ۙpA@~ �A��{�)bB���s�$$ ē~��,�kY��S@U,�f�J��(�JIzFId�����f�mf�h��3���*�`��v���hnzb����]�˞��!M�E�h7Rs�0=�U��9�<�*���L��0���B�DJ$q� Ɓ���(x� 2��]��J-����\�B0�7�3��b�� � ��X}��d ��Sg.����i��P؜G&��W�����@a�"���9*�Vn� CQ��j`�#C|���iD�H�������.]��Y5�C48���A���Yg��G�F6����O��&7ʙ� Z}���� Ҙ�L�Y2�H*  ?,r�a*���U��
Rbn��m�q�� ����wy�jĮԔ���&��G���SpU����i\��$�Aq&����e�����>z�ᴖv_�ޤԶU�}��������������tZ�T4���h ,R���)�&���"g�#��m<��#�/���L���N��B_�D;-^�~
,>��ۚ~OG���>�-fb;��M�K�I�
|o�A~T�7r$�����?��J��n�$�C�� ������K�FZs=z�>?�c��bpJ�4�x���b�b��N�J�����{�g�ٟ�p��f�Ѿm��D���*C���w��DQ�J>����D�qqbg������ke��k�gC��yV'�${b�9��'Z���CW�2&b!���X�!D�5M5�0WT��O�'ר�rz6�������z%���v!&,��ރ.sn����J=m;~I����3"��1kS{�ٴ3��	�\�^����Pω�^�@7=��×*=8�{����?5�>{�^�����Ǒ��)�+��G�����rQAAi^̳s� �`zc��;,4
�ۺ���q ���w��@0�?� Q����G��=`��{Q ~�|�r��ӓ|>�@��B���ߝXlE�] 6�!��$DSQ����ݨ�b(5-ǭ�ٽM+�tƟ�y���4��I�Pz|K[�I��@7-���}�Qic헆�����r�\�ָ_gQ�����5�2�^�ozS[#�;'�2��`���d#�M��+B�!��䙘�b}��8�e��I��U���#͈E���q��0{�3�~W��p!pl~�|�C/��t'{�}x�Q,Lt�aѠ��D�=i�Bl@)�}H��/ ~��ڒb�Ba|�^O�Ϙ8{T�fu�3i@r�Yr�B���zuҍ���Y�l�>Z�����|�?[�H06�(:ʠԠ���Q�-6��������V��B�I��Ǵ3�M8�k�F9�^8 �1"n��������-�'���O�0���,_p֓���1��s�D^��z��l���|j�:�s�܎���w�]�����c7E ��^!`Ƣ^ �������=@L��w�9�E���C�?��H7Eh�r���@�x��Ṽ;����B����6d�E*gY؅�@�����3r$kkb�bY���|�6��骭�s�t�D�� ��f${T�yk�j�E��(K]���3��1>nO�$���Mf*�#�Z|��_�2}l�V�I��1ɹ5g�x�D�܅�9Bxo�6�,(��{��
��7((��J%^ �`�]��P� ".D>��
�������ͫ�"^R�V�Z��_�$A:x~�Nr���
� ��+f҃,��`�z�w���3�샔���JO�
Q�f{�&ڹ'�¹����2Ϭ��n��'Ǒ��)��ޛ�yeâ�;�����O�͙~c�PK;���ͬd@X
�@�~�D����LW'Zf�>g�VM��3�xin*[�
KـU�`��f�̸�^{�&&n��*��JJ��f4ԉx����i�]�(��E�J:����$vDWiG,6g�[���O: \�R@�����ae`�$�X��0p\#_/`Ta�=AJ<�vn�7A�u���x\!@�X�P��?�9�܁w�K9E��p��7��
�q���s]���J�^{�|$�n}��Jy�.� P�*�0*���7�Ѿૹss�̝f�Xm��&�
��d*����~,�������g>y3������{+Xщ'��E���RkR�9�@�&2��c�t,.>c�E��|jЕ%��#b�K�}�H�^�5���¬pl~��}�=��$b����4  ����1O��;%�єG��HN-��2�P�����^�����V�W��\.� ��E�cck�@U&��NmU�{rv����8��9sF�u*����&i�;�FM/�3�b�w���)l<�3���K�[�.,J������zZ�
��>��]ѕ�����E����h $ ?D�ZX�L`nH��]��;>_�������L\Ĵ&!pOӣhN���� 0��L��ҋ�����]��m�/�=Dצ��v,�T��PG�������`�I>�W�v��i���ǆ:�m��W�V�����mi�]I����ޚz��h�:׋�9� :���h��U��و/�5ń#X3H_
�q0�a #!�s����G��h���C<����E|�U"���m�_&���h��4��6��'���@?zw�V���v`����7���<��C��N���Q�n�JJ����S�=b�33���hۇs�HkhR����N\*r���ҷ#��D���p����oL��^�o��~Lt���C��/�&�e����s"��dS9G�I�\��o xV5���0)E���0���/�n�T��NBH{�Ut�B��w�e  ��_��>��gD��PP�,����!t�	�� g�Of�@�}k3�؊0�`??�Xx��,��z�J��0�T��$%%:�7s��cFJ1Ĉ�ֽ�ԅ���i!�t�(zv�Z�]۩nDQ!hz�]��L=#�?>�d냋;�'��yS��[>_��*�n� )�Sy*�ekCD�Y5�c��§�|z��?���{:����N�+��w�5(v8)CFL�1�H�$mUN~�����B�����=�C+3�S��	T�7����CY~��ӕ7_Ꮳ@�����s�v,rw�:�}�^j:�{�+��׀� ��	�uN�+�@@H��"��,�0�Q�����	vu)���a-c��d��P VY}�ҡm��x �մ�_�Fђ�Fz>����2�i���t����rrǉ���?3~0i%�N�r+vs�>���h���r�33�Z�т�/�їf��g��u�����8��h�Ѧ�jV�`��	��b�����E�F*��R@��I�j��n�дr	'��TQYD~�u��/��C�ZZQN~EGxg��E<q�D��Q r�m��n��zz��+�W�0ʗ_��`Y�R@�yy�Op��$"��HM(c�	���Us�!�����=xI8a���B��-N�rD���>���TN�
��SCjMM���5�q�B���ChW�M�0Z��:KH��$z1�r����� �TI���4*Q�Ԍ�j9OΥzĶT5���	n��Qt�b���$V�u`q2d��|J~F�=\Y΀sr%h�7�	,�cRF�a��}�D`)`�a���)�X"��0z���A O�/\�
��3)[X.�v�P�@��[�3!�ɉ���ϓ^NwS��T(R��1�3խ*����P���wl�Տ[Nbpʫ�hD-v�[7ʈ����J�n���!��Q�����������U���g[��'JOg�&��(�Udè�`���! �AR"���� yL�4�"]M`PÀE���{�L��K��}O,�4wm�	�,);B�I/, Ѹ"CX��H)������m,�Џ� E�@��`�ɨ�*�競��W��k�>.�B.�Q9̃~X5�>t=�n��
�ʦ�cS&O��%��>�����#Z���HC=���Ϻ�`��'.Q�'�s9u��`�4qb���6����(i6�k+*��H[b�?��ڪ������?�0p��LqѸ� CD��Q��pX(R`���հ�p��x/��; �`T���x\��$�Q�wI
�� �� x_[��Z����X��F
�}�Ny��9_ʱ�S���Ʒ-��h��j}�G1�<YI���
u���Og׶F���C���Hf ��OG��4PR�4B'X�X���ҩǂ��g�f���Bb��7�7X
��ٗWy/O�|�|��w�C�j2Up&l���#���RzX4�1�4b ,jXRk���� )D^�����'�f#� wC��񡦄�E��o�����>�k�۩V� !ݗ�}�q����MXq��iF+�|?�Fˮ$�>�5!�����#�Eu��`�[ڛ(��D���9�t�m[BR��<��?��(��J]j&*������A~3NS��j�V7�؅����v�=�˞��^���,n,2oγ>���n�9p�}��@>؉���ɽ�>3�"XC|� �X6��׌�.��L�6�@41�)Dg!�ZA%z�����\iӔ ����
�y��TFб��}��꣄���ŋ�z���g  ���ݷ�j����[@���b燻�vR
�o��}Cay�ر�"A��!DO�wP�k�`�^G����{�D���6���!�����ͪ���@�M���� P������hz�1B]�kP���,QC�)�<s�f��ׯ��@lG�*�s� 1��� OaQ��,��ZJ�c�mȀ0��mg$��hCB���a��TYe���/�nl�H2��!�"�CIϙn]}T�ko23e4,��#���'�a$��e������7�J�&&n���G.eRKB�#W�������#k4�W'��3Qňb#��+1!8�vm����	�TPX�ݪӨ�:D�Ŕ�FU�njxD�"��5Z*k�	yJ�z��
��Z��몄�	R6�@i���/
e�D�	(9f�nmJ�x&��&bLpQg i3�2�Y՜�;���K��D��V���F�@�q}!%-�nЅ�|5L1-�����Qgpk{#�G�eɹ�u9���3@A��N�4�A�g�SV�ђ7.:t|u�g�XXE"�J+�Ձ���AY�Ӫ���ܣ�ʐ!���bO!�l�JEe�/�ᯱ�#��>��Ba�2���5g4.K�>��L�.���j�d�1В#Z�J��/��K�(4��.r���?ӂ��Sbt(��I���#5YD{˽X#C�(��*(l�X��4P��������.F&k���!�d0���c"�щc����欴f%�A}�Az~	���Wzm�M���)�YPJ�|��^��F���7�$���1i� 
�������0�[�/�#����y���B�]M0{�4z<!!ƴ5Qv��gIla�����,�B��0R����#����A�M�T2��}��B8����}F%����Y���O���S�d�L4t4F�3%e{t�[/�e��Q%�dp=3��N"�q&�vy���Ě�]��>n���֪H[�5Il��s�O�H�N��c�PCz���h���?X��C/�0�C�᫘@�M'^�
t>JEiU�VV㏕V��U����ۋoҧ�Y���~m�#�f��3���@����~��	F�㒭��@Z�e]"D���ƭW��lY�v�����{��^x��ZiH���Na6.Z�l�PӚ<�k��8�[��̰nm�DJ��"�F���V3S��L�#FT�,-����7Q�YM���hT�h��e\@�pӑBJ��(��n�H!A��!��~;�K�%�Ӵ����~���a�V��f�S[�y"5��������=0-Td��`kvU���s���;�Ƙ��Q��｢��� o�I+�8���gO<���^��/�|%�߸@x?��&�Lg�\����ߏ���z'�M7�Sk:u9����ؙz��a#��}aM1t1�(��Ml;YD���Vd�V/������#��~.����|��Lٖ�M�"�'ﭠ�����VQz�
�dvޓ@߽:�5�A�G ���b#)�
&��G�|�V�@L��dA���΃�?-�X:w���מ��#�l���.G_��FՁBD�P9N�1���Dop���+����-�JP�BL�酫k�&`��~/��M˶u97�Ǯ�D��XNM����Y<�8�O��%��L/CF�|�l�	J!�{&�n�S'˞�^�A�B�v��n}m�M�k�֣��d�E��֑!t.�u=�����2e��E��G.�7)>���!&X�.��G�����o���B���ݷ�<o�4g��:���"�����V�ßv�'��/�4P�������r�K2@��7:�2�}�U����vsJ*��-�����*��J0������@|m*�j���.���`w �R�A~�ḅ3{��t�S�'�|.�O��Bv����^�D1a�Yd0w����(*pX��肝�_�QL���H ӎ _&��CRL ��-e�V�˥ml iҌd�:O�c�uI��;O���Nӎ�VT�\���,&D�H=Hk�t����E�1��p�9�An�c`�̈́H���8���ʭ�"���J ���`Z��U�啬�@?��f�i-}�>z��e�_�=B�4��-[��DR���t�P��RM�XDj��j�!r��7�Dp��\�2�wE�К��L"]I�B��Nn

�3hEJ+��)��'Sh��34��;�a�CaPq��ا�QJ�{��i7��ߢ��f�~�����.�O�=W��/�ۮu2H/U�1N��I�����3f��`����Gf͜�5�x����^�R�>j?��B"���7���G���y|,E��<�&���� ��1��V��ё�_��\��� �h�U� #��O�L��rQ�%K��>6�G�N����2��������E����x&m,h�𸑳�}���ð������㟥�L�S�D��!c6(��/ô�;�-����5O�<ci�P�É�)P��d�2��*V�$2cژߍ}��rKs�:���O�����!�5�/C-�a��l�Nf��)C�	�e�ˮ��\�v	�&�Ǔ�h���	P��0��m|��N��� �*.���r�b��PX�`���mWq��U5:��5����%���ǜ�gQ�n`y�C�I4�!6\H��hs����BB�hs_��o�����D��H��p� ''�����!�jĺ���w(
В�8#��q^�|�H�:�!JU�B������G/YyXPĲd-UzX���s���
�&8��_Ia�~zqY��a2Z6ΜO������כ#�uH����4t[{/e�X�6*��WҪ�Z����#B�Z����N�J��;|!�6��t�����N��R񢣂�
�T4� �'PI����5��5R���v��.�Y��'Í �gG�L�H.��f���J�=�������gx*pr)��}oɐ!�=�5Í�J4���t$�0��Ή p{,�w���f���D��,6�L��^����*�}E��l	hצuL�>����K��"UL�z��|����`�3��4jxw����+��Gλ|�M#z�V+MO�7���G���D�ҧ(���ۭ��SR�m-�x�����e=����&�L4S�h���E��En�b]�U�;�Im,�i*vCP1ԗ"1���]���1�&�q���c��"�Vѡt��!$�7pM>��w<9�-�q� 
�6�����-��+u� �w�=��uI����%������� @�~�y5���7��J���J�M�Bx���7/g���M �&��r=�`�S,-�� ]��-��D�.�*��
P̣h��f�&��� JD��7����7o�//�.8 �aω,Z���Ρb-�{�
�K�H��w65�V��B�x:���F�Ӱ�1�-��J�ۣ
�b�d��ҝ7��d**��2:m�e.bW��40�����9��,�L��e6=�GI�a�-�ˢYqdP�q�bM�XJI�$C�
%�C�Kt�%�2��j�2ڐ�fa)��:�Q�Udiy}q6���Uo�я9�U��b�|~",�/��)�R],cR�h{Y;
=v�F��`V,�S�����y�КVH��{���h6�*���L�Dӗ�r�1�Τ��O9m��I��BK�h�=����fR���f-�ֿ����ӗY�aܠ.��>ɩ�t���1���}-�0���\.�A�<'�sW���!=�2x~~9�e8.���~4���1r9�o�pre;Oo��E�@�5����R�S�0;�*9�ܕ��Iz��z�UA�/�������=���U���p�����6ѷ����^�y8YM�']}��C���f?�U�G��e�RJQ�s��;�OO�y�����w�se!�Ϲ\���ǳ���ϭ0��j�Zk�SP�vy<`��b����V���A��5����񶧩8B���f���h%�jj��F�����
*��<�*�U�v�s$�W�C�s�ؙJ�e�W;$��}Z��S���|�,��`"�O��H��r˽�Io�ۑ�kK�5{N�J��$����������z�6�x�ڑ:���� .�l7�T)�V��?���5.� P+����r(�r*j.0��и�[$����=��S��x�a�컐��p�WѦ�ww�c�ܜ�q#w��.�;���"����xͱt��qi�vj}��d=��L		��=�AN��N�*�ڔ��sKH!��`b�����xc�p2��3��5�;�f$�	����D �@��8Z�����9�iT�ˡː���oaC��� 	��Vo�c;is���HQ�n�����x�K�hQ�31v�"rf��V��&]�ˁ3TRQש�����2�a�h�4apW6L��ʴ?�u�C�H=�C����A/CR���8��
��������]s������^-�Kƚ�S�DK�9�z~��t%��Vl;�ì���Ay%�T$7ɸ��!>��=�v2 ��D���2<,��܄Gz�I��&�����z�p�E�wQ2�{L�m�x �0�����I�38x.�^\���}b,�q�kJ�1��Q�G��-U�`d���2���w��ߗ/�Ok��#�ӗs%�զzA<⃬4�s-��`Q2�cf=b�.W2J�;��%���:>��G�[
�-�qLt0SZ����ٌ�T�2�wWm�y?lc��d�h)��=����{�AZ��4�O$�������DVS�UŹ��l�\nC��&�:�~�
0�s�w��ؘ5!DW�D�^�}�}[��G�߰�6�7j�uײ�����7�?T�Y�h�4~PWҨ�ԯC��4�$��;�VU��km�B)28�_H�t��;q9{@�pk��<+���^�H2jbn-��=�O\uʶ��a�"
�h�'�җ�� �:6n�3Ǵ�#�Y�O?�1�b����F�!*]�4}�☋ V.;et?��\P�~�W#07Ag��)>�>��D:r1���[�jiܡK���"a����W,�����n��ó�t��D�[l*�E���S��ف�-��������c.�N�p�m?܍�J�!�]'S���9��tiE�L��V��!z�?�Zd�hn`���D��=���FW)��q�ˌd=�a���5_}5���W�/����鈂}�6�Md�u\�HE�m��Չ.��pO����~�!�KÙ�d���˺�ͯ�[Χ��os~�"�)�dʐ��8v)����tۍ��9�[�_�(($��r�E��L��y���tn�@A$'+$=O�}��*,���|h��˜)��Sd�h(9�Bo������t٣K5��D����lzI�Ud-I�D5������9ȠXt�ѸȄI?}�����?���(�Kˁ��HeW�ؿC<}<�nF�s~��Z?b�!���I� 4`�Bf�~���,F����a؊;�T9Q���~|f����w"Ԏ�q���٭M2�\��F�az���Y��D�������8�����$Z1`��݄Z2�F�%�j���y�v8|��oY'.&*}��D6�}���:W�\*�Q���.a���L;�8cFHb��	����ܐ,BB���n�~:���iӆ�]X磌zt�O���?ڇ9Υ�t�B	�v��,���v��-G/�D �E 6,�sα�9�~�I߾� ���%��y*V9h?���y���_5o��$�˧<7;�uh��p?����	MDј��T5M��ز֧��{b�2�k�鍊>J�,��k���:DAẠ��>���iߙ��SA7tN��}��xJ���52�%��n(g��4�3B8a�e5�L��Q�8<�4�ݿ�ݕS��ùy���&������`��Yi{��!*�rTt�P�j���cQ���@�ǁ�NS[��H�2|��ެM�˹E�ˁ���۫��Y�����vʐq-"�OG��z�5-=u� Z��Vl�̄���-,�VG��	����Z��M7�;��P�D��D� �×Ǵ��z
��?W�:�!��>L���~����}��݌��C����z����\�(㚂�fj�������o�� x�:ĳ�X^�42@�]��-@rl���y8Q�Ԡ������z��,�w�Ԗb��N
L��E�Ʒ�1=��7�Y�����=������)F�d\K�q���d-�x\�-f�~��A�a�q�MJ<0e�a-s��<�>����Oh�<1��3�������^�!�&�L� u�傆�������C;�SH��k��a�	��Ъ�-��h�^��h��f������vr��ž��{�mMUS�h3����b�+��G��q�g�$eĐST=4��;�ѿ��Nێ_b7 E��:�YeU�!CF5���Q-�X�G����`m��e�S�������U�a�� Yy�m!���@-��+6����H��_��;^{`4�hӊ5s�U6���*2ʔ춱���W�:2���{�DJ6K#
�t���Ct2-�dȐ�xP+��ܫe������2���y�QB�T�g��ɐ!㚆^�&�W�V���}��Ƭ�m!��`*�2dȸ�`Q(�c�k�]�$z6p�sȢz���Y��O��!C�5� b���࠿C�O[���J�׈�I�-�ل�%D_Ҝ9_(��)Xiɐ!���ujq�K)�Z��g#�e6��D$�8�!��Ar�A��wvp���0���B�8kag-xP-C�����4sϦ��:c�Z�}ʪ���H!�dȐqM��
Ċ� .0'��i�L*��V����cI��$�]�\��I��O��|�_�g����~�(�.C���כ�eN�
ƿ�Aa�i$C��k
ި���9� CƵ���ZTpv��dȸ�pմ0_�����@+�,��d��� R�Y��J��cniUV��P��d%��J��ʸs�(Q:�ՒquC&�� C�Mtk���5�����Դ欆*�QR�"��H��̤�@��*MD\����l^c�ɠ�1����'��T*��ǚ(!�L��4!h8k��~��:��宨;8�,�oNhI��w�@&�fD�p���&:y6����%�Qtd`�cQ�V�����%7}���LD�_XA�.�F�����߯n�N�Vf:�g����%v�@�K5#���%��L߯;N�eU���2趛�PB\H�s��2яg�MCPq��q�?�sKi�Ɠd��p�t&�;�������f��!��fD|��}1-�� ���NfؐfL��.6��Z��.�q�tV- �dΜϥ>=�&�s�Bu�QƵ ��
�eb��O�ĉ���Z����k24#2�T��3�۶�G.SeU]��k�h��`�e�5-TK"�ȣs�h���_ DܠC���e�+d���L͈=�*D��뫡���`���j���F>�)a�`���@y���c�ҙ9��w���@���{ӛ���έ��>��<�ΧK>�'�kFɩ����A���l�`}�-�]�̣*�g��d2hF�Q�!n�a�.�� �V��d���摐�pNCB�,��#�#��p&OE{�4����_嵐]۸|�'���[��p{,���f�$6�g��ElRxC����1�qw2��t]���B��x�}.~V�T�dЌ���,YK��F�h&�ʹQ�ŵ�ƣ��	}�_G�bdc����w��i�y5w!�Wǝ��>Y�W��:�Sc���\���&Q϶�����IC�W�a�U�o��}q1��X243�`6]�����v�_b�{f+X�+(�X���570���cZ
�RB��"��� 
�(�\s+��R�l�*I{��6�O_�v��{e2#�
�������z��!��D:M�/g�[������2\%Л�Gf_��RTum��+d������6���=����='��`��G�j��(*���此����v>#��^�8'=�C&�5@�U���i?^H3��>rK����G�7ر���=A����9�$�*��bC�+W𥏧�E>Zv��g��y2�f�;��"�����J}����X���C�r�����#��}�q���
;��M���&��v-sXĽotH ���5;��C�<��MF�"�42�D��Rqd�[���jښ�b�+2�&l<x�2�Kh��%�!.�wI�|w����Hn�������K�BBT(��c�Ș>I6dгm+��!���&�҄Zn��hÈ����a��Ǌd��Q=�7�y#�<јq&Fk;�i|G#�J�hD�Y��$#��6�'�;�p�ث}��&��>^�����~��ى4n`���9�F����y�-��I7�/8��RS筠��*����x�f�C���W�PRl8}�ܟ�
���9K�̕\��2�ˁ3��-��z�.p���ˮ3L��[̮�O�IO,XŞ7�_P������R�{���xC]F�O��/_�D���D��r���F>7��)uK�fiJo �`{�&���w
� �k< ����ZE�V���@+���@�qL״����o��.!2��MJf�����?v)��Nۼ�̕�@�����'���{O�ɴlR+U,r�5�E����,'֟��V�׃�K{�Ùy ����������|�}�9�$C�+|��(�=�;��9�����]S��?C}��'"��sʻ���gP��q�Pht7��v�[>���ͧ)�J�"B���[�Qp�u�\4�d�����I����w�Sw��� 8u9��q!�<X	�?����~�����7�j2 &���畔ӧ���{���� ?�ϕ!CU��뿤�������Կp��н �J�Z+E�T��\.�%������G���~G�=������q��&)�9ߞ3�T��X�%���ߒ2lѨd���ܱ�Tp���3	����>��<�b^]���_ʬ}l�׿�w�N�u���_��;u9�^[�Km�,�xg�V�~�ɐq=�Qɠ�[�&�&��:v�r����>��J�B�v1�����Z��q���*:��ͽ����m^{1���{�z���9(��אn,
���?��9S�G�jv�� ������S6yS�$�[ChN��6���;��<���;V��'F�D�Z_���h����2L�UQ�h3�����%�k`0��}�p�ս�KЛ�N;��Cj7�����2������ESE�����<w��y|,u��n�5MN_/�eD��~���-5*jR�|갂����˄�8_߄��g&�� ����MQ������~�A��P,UY������g�$e��{�����O`�3�MU�@\NM���h��n�����5᳍����F�u�yO���mZ�/�B�����b�&ű4�%�J�Տ#X�N�`-Xp=j���̸�t��N,c5�6�!W߶��GX��7��HT���+3����)Y�����Ѕ�r�׿��m`�kۉa��j�i�c#��Ug!�ɩ��m�/��w�q������렜����ϯ(&�N3���ң��F'��J%-:��G{(���\�����v]v~���� \�������Nz|�*��5qp7��_'��`�Ga�?�����2�6��8�c�� }u�/��SĢ�����3m^�/��~ɊNj���R��l�k�Ǆ� "���wl1	��z�c`g�������\���%���<�R�s.��
�WlJB�<p?C
9�}��'�bh�
�+%Jz{���2S�`S��*W��lkzq�7��A��u����B��o���hP���%�V����?��>�UWT|a��e?��i�������>��uۺ*�q�R�a��:}i�O��@��d���A-MV��@��,�I�X9��I7��n��]T�JJ�p%������\h��	�U]���t�]O��eȐ� ��2d2�!C�L2�L�s(��%�zg9��;҉&A�`��x�G�d � dϟ�0��K�%�b��!]����)�p�&%�ZD�Y؈0|�=�l����0��j��_X����C>+��X�\#��m�t)t-�e��z<���в��������m�h2 	�nk�	&�ه��x��֞ո�5h	 	�7�� XW���(��+�'��g�7��qCf�A{:���/����G��#RP)�4iT/&H�l�I��}*�Vl?�L�ރ��,�u�3�@��6P�[f��;�L�C-��喷\B�����ښA�^:GX�m��Uh��B���g��)@k���;ԭ�ʹ��N2!�ܚs�iŶc���y,�a�5�;�u�`Z��x�^�;$F�Ҕ�}飵����������(�OG_�~�Z"��{����k4��M�P
�c�����}:j�վ�b�D �NE4���Uh��K�]� �O��HBt���p�Jܚ*���;��k�h�%���4id/ճ�dM�q;���!]۰� �]C���'�12����<� ���8W���Bw��B1�A�:��ʔ/��ݑǈD����0��d_��`�A��F��N=�Ų���3�=>�U�� 2@{�T2�[tM��of?@�n��z��P*Z�ۨd����|1%�� L�9r"����� �@\`�v_ZVE���3�'Tńe^��]��E�Ab��ys�b.��C�O�8f!�V
䮍R	��:�G�>�w@/:
�u��Q@���Զ�C��M}0�� �\�^B�L#�VD@s�]#��&���T!�;랑L�\���R�ײ?X{��~?�a�g��i�M ��A���#j%�x�LNaZ���Q�@���!�"6��>U$\������_��������^Dz������jh��2|$��8y6���X�{���Ћ�jfj$p?��1)���HNɦ�������d�O���0���~i�gh5�V�@���};П�������׶CsɌ{X�������,��1	�[�ڪ�p7���������f����  �Z�1NHD<pnWWU�!�6!��Nc��G����?g��<6�Z�>SzVq-�8s!���ʖAje���`�b�K�\�,"�����&ڈ�o�i���9����D�jS���v���݆���Ғ���~eb% �ԗ� ��t����'�adЛso@X��D�H���r����&�Ĉ�M�r��`�����)*c?C�D���,��9�5���J��{ KMC�MLy�m��0�` DR��خ��Z<Wز\@x���f 4��Z u(�|u�ՙ�R>3bM0�c�b�O��ߋV&*�u礭9���ǿ?bs^���"���{"��R�fWB'��rn����X���Z� �3���Z�VB8+����_�;Yr��;H%li��<Qz����yu
�P����B�h��6�ǂYqR�"�*��=4 �#�� �]�u&���`�ٻ���(#��V�;4ؗY�<����5���h;��݌�Ӂ��E[��Ǆ3�H��@p�����y�mH`A�X�-�˄Z2��Go�Ojn�C�q�o�K>Z%�f3��� �����D���r_���r���~M�j�Nv���[�����~�L&�����x?�D���C�J������禗���c@�@yF�w�ѓR�
��G��B��Z�4Jc��ú��Gn��Lg{�S���Ӂ`JÜ?~)���e�51��"6���K惙0ב�@�c�q̧�(�x���k��@���{Ӽ�Q��x����,�~�~@eUՃ`��}�S렬��Ａ+��I�&�@,�->�e3�BԨ9��LI��dn�ug�~x�PEê��cg�rK!����Y���#�#��ؘ?���!4���L�J�{"��M}�Ϸ�L�~;�2��V���y���LC��Y�"�لi�]C��U�1�+7�C��h�8�>{��~QX$?�1�V�,��#ơ�G|��u����큛�M���.Ҕ��ђ_���A]��2nB@�.��h�ބ�rwk�T�zQM82p��p�x��eXɟ�U��	W�tQ�������k�Y������"�Xѡ���7�!98�ᖾh�˓�X3� X,��q�w%�ca�����Ɣ[�[BT��f�KL���>���ə�H��9Ag�Go���"�&��n�����8�+��t���s�o9B˹�G���u2�Mm�Q��x!3���b|�o�kAR�kΩ����������?з.�����F��B%�>���:E	!�BA_׶���ҷ���?�F���x�)`�<���O����n by�4�hn�����Y)1����M��6�47A�|���;}/L�b��v@��p;�U����v~T0�t:�&|��~�
�Ґ��d2h켬f��hTJ
5s� QA��e�iK���uo���p�K0Q�X3E�YX���"mIQy��F�������fh`��tTb�y�v1,;�����@�k�d�DH-V�gG�ue#��7��٭!3>�&'������2Ȑ!�A&2d0�d C��dȐ� ��2d2��V���
�e�R�u(l�:�ia�~s�F��`0z�J�B�7�6�|����7��|�M+�߹_��&�L����V�v�\g���E�F�Q�j�^�ԑt>���.t�`&�>�� ��nY���&�L��Ii�N���Q�^`�B�bܬ�9�]L2�2��c����d���C��@�+������$?_a�k��l�j!�A�'���<�������������L����򸐐�Z2 ___���X&S����ucǎՓ��NV��R��m����{FFFw�=����AAA��fs ]��j�`RO���~�w����$�@���Ym٩6__��ؼy�����3�Ѹ?<<��ွ{�NT�T���O�'L���d47�N�k�]����Qt��s^��-w�#����8*%??��<��x�U$��`���3���
R�$���_�������;�d��_�~k<�����~�<����7��l�*hn��A��s��{i�����b�Z�Ӹ|1�"�>dȐ�7u�
�Q�w�m�v���j�����;V"h�.�����M(��|`eb(�g�Z"d��p�������dHƈ#~���Q�1�U�mU�[���ևK#fP��+��L	?k�ªx��'�Z���=m���ˮ.��ρ�q��j�J��zTA�wK~�Ϸ�5BЍ^gP�v�'t��/�T�(,�V�5��uXgK,���FG��s��O�5��-k3i.(IUa6�/Ul\�0l���.��    IEND�B`�PK 
     T\:�b��N  �N                   cirkitFile.jsonPK 
     T\                        �N  jsons/PK 
     T\�#��(  (               �N  jsons/user_defined.jsonPK 
     T\                        <_  images/PK 
     T\ѥ� �� �� /             a_  images/41d41cfa-55db-4eb2-805f-824b346b9186.pngPK 
     T\�j�ؖ  �  /             E� images/2dd0ce04-414d-4887-acda-26c206c9abda.pngPK 
     T\,b��9F 9F /             (� images/1d10c801-e2f1-4174-9a9c-587482dea60d.pngPK 
     T\�,9__�  _�  /             �= images/05c4396c-27e7-4cac-a4cc-0e5db7270844.pngPK 
     T\��v�z�  z�  /             Z� images/f814d8c7-8d80-4469-af20-bcf736e1bcac.pngPK 
     T\��  �  /             !� images/858a2a89-b1fb-4d30-9067-568b89f7eae7.pngPK    
 
   �G   